MACRO cell_0
	SIZE 100 BY 100 ;
	PIN pin_0
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 89.68027888446215 0.25 89.93027888446215 ;
		END PORT
	END pin_0
	PIN pin_1
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 89.36055776892431 0.25 89.61055776892431 ;
		END PORT
	END pin_1
	PIN pin_2
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 89.04083665338646 0.25 89.29083665338646 ;
		END PORT
	END pin_2
	PIN pin_3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 88.72111553784862 0.25 88.97111553784862 ;
		END PORT
	END pin_3
	PIN pin_4
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 88.40139442231077 0.25 88.65139442231077 ;
		END PORT
	END pin_4
	PIN pin_5
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 88.08167330677293 0.25 88.33167330677293 ;
		END PORT
	END pin_5
	PIN pin_6
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 87.76195219123508 0.25 88.01195219123508 ;
		END PORT
	END pin_6
	PIN pin_7
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 87.44223107569724 0.25 87.69223107569724 ;
		END PORT
	END pin_7
	PIN pin_8
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 87.12250996015939 0.25 87.37250996015939 ;
		END PORT
	END pin_8
	PIN pin_9
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 86.80278884462155 0.25 87.05278884462155 ;
		END PORT
	END pin_9
	PIN pin_10
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 86.4830677290837 0.25 86.7330677290837 ;
		END PORT
	END pin_10
	PIN pin_11
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 86.16334661354585 0.25 86.41334661354585 ;
		END PORT
	END pin_11
	PIN pin_12
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 85.84362549800801 0.25 86.09362549800801 ;
		END PORT
	END pin_12
	PIN pin_13
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 85.52390438247016 0.25 85.77390438247016 ;
		END PORT
	END pin_13
	PIN pin_14
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 85.20418326693232 0.25 85.45418326693232 ;
		END PORT
	END pin_14
	PIN pin_15
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 84.88446215139447 0.25 85.13446215139447 ;
		END PORT
	END pin_15
	PIN pin_16
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 84.56474103585663 0.25 84.81474103585663 ;
		END PORT
	END pin_16
	PIN pin_17
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 84.24501992031878 0.25 84.49501992031878 ;
		END PORT
	END pin_17
	PIN pin_18
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 83.92529880478094 0.25 84.17529880478094 ;
		END PORT
	END pin_18
	PIN pin_19
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 83.60557768924309 0.25 83.85557768924309 ;
		END PORT
	END pin_19
	PIN pin_20
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 83.28585657370525 0.25 83.53585657370525 ;
		END PORT
	END pin_20
	PIN pin_21
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 82.9661354581674 0.25 83.2161354581674 ;
		END PORT
	END pin_21
	PIN pin_22
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 82.64641434262955 0.25 82.89641434262955 ;
		END PORT
	END pin_22
	PIN pin_23
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 82.32669322709171 0.25 82.57669322709171 ;
		END PORT
	END pin_23
	PIN pin_24
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 82.00697211155386 0.25 82.25697211155386 ;
		END PORT
	END pin_24
	PIN pin_25
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 81.68725099601602 0.25 81.93725099601602 ;
		END PORT
	END pin_25
	PIN pin_26
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 81.36752988047817 0.25 81.61752988047817 ;
		END PORT
	END pin_26
	PIN pin_27
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 81.04780876494033 0.25 81.29780876494033 ;
		END PORT
	END pin_27
	PIN pin_28
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 80.72808764940248 0.25 80.97808764940248 ;
		END PORT
	END pin_28
	PIN pin_29
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 80.40836653386464 0.25 80.65836653386464 ;
		END PORT
	END pin_29
	PIN pin_30
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 80.08864541832679 0.25 80.33864541832679 ;
		END PORT
	END pin_30
	PIN pin_31
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 79.76892430278895 0.25 80.01892430278895 ;
		END PORT
	END pin_31
	PIN pin_32
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 79.4492031872511 0.25 79.6992031872511 ;
		END PORT
	END pin_32
	PIN pin_33
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 79.12948207171326 0.25 79.37948207171326 ;
		END PORT
	END pin_33
	PIN pin_34
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 78.80976095617541 0.25 79.05976095617541 ;
		END PORT
	END pin_34
	PIN pin_35
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 78.49003984063756 0.25 78.74003984063756 ;
		END PORT
	END pin_35
	PIN pin_36
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 78.17031872509972 0.25 78.42031872509972 ;
		END PORT
	END pin_36
	PIN pin_37
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 77.85059760956187 0.25 78.10059760956187 ;
		END PORT
	END pin_37
	PIN pin_38
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 77.53087649402403 0.25 77.78087649402403 ;
		END PORT
	END pin_38
	PIN pin_39
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 77.21115537848618 0.25 77.46115537848618 ;
		END PORT
	END pin_39
	PIN pin_40
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 76.89143426294834 0.25 77.14143426294834 ;
		END PORT
	END pin_40
	PIN pin_41
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 76.57171314741049 0.25 76.82171314741049 ;
		END PORT
	END pin_41
	PIN pin_42
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 76.25199203187265 0.25 76.50199203187265 ;
		END PORT
	END pin_42
	PIN pin_43
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 75.9322709163348 0.25 76.1822709163348 ;
		END PORT
	END pin_43
	PIN pin_44
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 75.61254980079696 0.25 75.86254980079696 ;
		END PORT
	END pin_44
	PIN pin_45
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 75.29282868525911 0.25 75.54282868525911 ;
		END PORT
	END pin_45
	PIN pin_46
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 74.97310756972126 0.25 75.22310756972126 ;
		END PORT
	END pin_46
	PIN pin_47
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 74.65338645418342 0.25 74.90338645418342 ;
		END PORT
	END pin_47
	PIN pin_48
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 74.33366533864557 0.25 74.58366533864557 ;
		END PORT
	END pin_48
	PIN pin_49
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 74.01394422310773 0.25 74.26394422310773 ;
		END PORT
	END pin_49
	PIN pin_50
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 73.69422310756988 0.25 73.94422310756988 ;
		END PORT
	END pin_50
	PIN pin_51
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 73.37450199203204 0.25 73.62450199203204 ;
		END PORT
	END pin_51
	PIN pin_52
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 73.05478087649419 0.25 73.30478087649419 ;
		END PORT
	END pin_52
	PIN pin_53
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 72.73505976095635 0.25 72.98505976095635 ;
		END PORT
	END pin_53
	PIN pin_54
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 72.4153386454185 0.25 72.6653386454185 ;
		END PORT
	END pin_54
	PIN pin_55
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 72.09561752988066 0.25 72.34561752988066 ;
		END PORT
	END pin_55
	PIN pin_56
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 71.77589641434281 0.25 72.02589641434281 ;
		END PORT
	END pin_56
	PIN pin_57
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 71.45617529880496 0.25 71.70617529880496 ;
		END PORT
	END pin_57
	PIN pin_58
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 71.13645418326712 0.25 71.38645418326712 ;
		END PORT
	END pin_58
	PIN pin_59
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 70.81673306772927 0.25 71.06673306772927 ;
		END PORT
	END pin_59
	PIN pin_60
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 70.49701195219143 0.25 70.74701195219143 ;
		END PORT
	END pin_60
	PIN pin_61
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 70.17729083665358 0.25 70.42729083665358 ;
		END PORT
	END pin_61
	PIN pin_62
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 69.85756972111574 0.25 70.10756972111574 ;
		END PORT
	END pin_62
	PIN pin_63
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 69.53784860557789 0.25 69.78784860557789 ;
		END PORT
	END pin_63
	PIN pin_64
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 69.21812749004005 0.25 69.46812749004005 ;
		END PORT
	END pin_64
	PIN pin_65
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 68.8984063745022 0.25 69.1484063745022 ;
		END PORT
	END pin_65
	PIN pin_66
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 68.57868525896436 0.25 68.82868525896436 ;
		END PORT
	END pin_66
	PIN pin_67
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 68.25896414342651 0.25 68.50896414342651 ;
		END PORT
	END pin_67
	PIN pin_68
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 67.93924302788866 0.25 68.18924302788866 ;
		END PORT
	END pin_68
	PIN pin_69
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 67.61952191235082 0.25 67.86952191235082 ;
		END PORT
	END pin_69
	PIN pin_70
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 67.29980079681297 0.25 67.54980079681297 ;
		END PORT
	END pin_70
	PIN pin_71
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 66.98007968127513 0.25 67.23007968127513 ;
		END PORT
	END pin_71
	PIN pin_72
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 66.66035856573728 0.25 66.91035856573728 ;
		END PORT
	END pin_72
	PIN pin_73
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 66.34063745019944 0.25 66.59063745019944 ;
		END PORT
	END pin_73
	PIN pin_74
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 66.02091633466159 0.25 66.27091633466159 ;
		END PORT
	END pin_74
	PIN pin_75
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 65.70119521912375 0.25 65.95119521912375 ;
		END PORT
	END pin_75
	PIN pin_76
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 65.3814741035859 0.25 65.6314741035859 ;
		END PORT
	END pin_76
	PIN pin_77
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 65.06175298804806 0.25 65.31175298804806 ;
		END PORT
	END pin_77
	PIN pin_78
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 64.74203187251021 0.25 64.99203187251021 ;
		END PORT
	END pin_78
	PIN pin_79
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 64.42231075697237 0.25 64.67231075697237 ;
		END PORT
	END pin_79
	PIN pin_80
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 64.10258964143452 0.25 64.35258964143452 ;
		END PORT
	END pin_80
	PIN pin_81
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 63.782868525896674 0.25 64.03286852589667 ;
		END PORT
	END pin_81
	PIN pin_82
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 63.46314741035883 0.25 63.71314741035883 ;
		END PORT
	END pin_82
	PIN pin_83
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 63.14342629482098 0.25 63.39342629482098 ;
		END PORT
	END pin_83
	PIN pin_84
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 62.82370517928314 0.25 63.07370517928314 ;
		END PORT
	END pin_84
	PIN pin_85
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 62.50398406374529 0.25 62.75398406374529 ;
		END PORT
	END pin_85
	PIN pin_86
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 62.18426294820745 0.25 62.43426294820745 ;
		END PORT
	END pin_86
	PIN pin_87
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 61.8645418326696 0.25 62.1145418326696 ;
		END PORT
	END pin_87
	PIN pin_88
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 61.544820717131756 0.25 61.794820717131756 ;
		END PORT
	END pin_88
	PIN pin_89
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 61.22509960159391 0.25 61.47509960159391 ;
		END PORT
	END pin_89
	PIN pin_90
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 60.905378486056065 0.25 61.155378486056065 ;
		END PORT
	END pin_90
	PIN pin_91
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 60.58565737051822 0.25 60.83565737051822 ;
		END PORT
	END pin_91
	PIN pin_92
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 60.265936254980375 0.25 60.515936254980375 ;
		END PORT
	END pin_92
	PIN pin_93
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 59.94621513944253 0.25 60.19621513944253 ;
		END PORT
	END pin_93
	PIN pin_94
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 59.626494023904684 0.25 59.876494023904684 ;
		END PORT
	END pin_94
	PIN pin_95
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 59.30677290836684 0.25 59.55677290836684 ;
		END PORT
	END pin_95
	PIN pin_96
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.98705179282899 0.25 59.23705179282899 ;
		END PORT
	END pin_96
	PIN pin_97
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 58.66733067729115 0.25 58.91733067729115 ;
		END PORT
	END pin_97
	PIN pin_98
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 58.3476095617533 0.25 58.5976095617533 ;
		END PORT
	END pin_98
	PIN pin_99
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 58.02788844621546 0.25 58.27788844621546 ;
		END PORT
	END pin_99
	PIN pin_100
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 57.70816733067761 0.25 57.95816733067761 ;
		END PORT
	END pin_100
	PIN pin_101
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 57.388446215139766 0.25 57.638446215139766 ;
		END PORT
	END pin_101
	PIN pin_102
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 57.06872509960192 0.25 57.31872509960192 ;
		END PORT
	END pin_102
	PIN pin_103
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 56.749003984064075 0.25 56.999003984064075 ;
		END PORT
	END pin_103
	PIN pin_104
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 56.42928286852623 0.25 56.67928286852623 ;
		END PORT
	END pin_104
	PIN pin_105
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 56.109561752988384 0.25 56.359561752988384 ;
		END PORT
	END pin_105
	PIN pin_106
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 55.78984063745054 0.25 56.03984063745054 ;
		END PORT
	END pin_106
	PIN pin_107
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 55.47011952191269 0.25 55.72011952191269 ;
		END PORT
	END pin_107
	PIN pin_108
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 55.15039840637485 0.25 55.40039840637485 ;
		END PORT
	END pin_108
	PIN pin_109
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 54.830677290837 0.25 55.080677290837 ;
		END PORT
	END pin_109
	PIN pin_110
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 54.51095617529916 0.25 54.76095617529916 ;
		END PORT
	END pin_110
	PIN pin_111
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 54.19123505976131 0.25 54.44123505976131 ;
		END PORT
	END pin_111
	PIN pin_112
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 53.871513944223466 0.25 54.121513944223466 ;
		END PORT
	END pin_112
	PIN pin_113
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 53.55179282868562 0.25 53.80179282868562 ;
		END PORT
	END pin_113
	PIN pin_114
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 53.232071713147775 0.25 53.482071713147775 ;
		END PORT
	END pin_114
	PIN pin_115
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 52.91235059760993 0.25 53.16235059760993 ;
		END PORT
	END pin_115
	PIN pin_116
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 52.592629482072084 0.25 52.842629482072084 ;
		END PORT
	END pin_116
	PIN pin_117
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 52.27290836653424 0.25 52.52290836653424 ;
		END PORT
	END pin_117
	PIN pin_118
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 51.95318725099639 0.25 52.20318725099639 ;
		END PORT
	END pin_118
	PIN pin_119
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 51.63346613545855 0.25 51.88346613545855 ;
		END PORT
	END pin_119
	PIN pin_120
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 51.3137450199207 0.25 51.5637450199207 ;
		END PORT
	END pin_120
	PIN pin_121
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 50.99402390438286 0.25 51.24402390438286 ;
		END PORT
	END pin_121
	PIN pin_122
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 50.67430278884501 0.25 50.92430278884501 ;
		END PORT
	END pin_122
	PIN pin_123
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 50.354581673307166 0.25 50.604581673307166 ;
		END PORT
	END pin_123
	PIN pin_124
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 50.03486055776932 0.25 50.28486055776932 ;
		END PORT
	END pin_124
	PIN pin_125
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 49.715139442231475 0.25 49.965139442231475 ;
		END PORT
	END pin_125
	PIN pin_126
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 49.39541832669363 0.25 49.64541832669363 ;
		END PORT
	END pin_126
	PIN pin_127
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 49.075697211155784 0.25 49.325697211155784 ;
		END PORT
	END pin_127
	PIN pin_128
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 48.75597609561794 0.25 49.00597609561794 ;
		END PORT
	END pin_128
	PIN pin_129
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 48.43625498008009 0.25 48.68625498008009 ;
		END PORT
	END pin_129
	PIN pin_130
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 48.11653386454225 0.25 48.36653386454225 ;
		END PORT
	END pin_130
	PIN pin_131
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 47.7968127490044 0.25 48.0468127490044 ;
		END PORT
	END pin_131
	PIN pin_132
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 47.47709163346656 0.25 47.72709163346656 ;
		END PORT
	END pin_132
	PIN pin_133
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 47.15737051792871 0.25 47.40737051792871 ;
		END PORT
	END pin_133
	PIN pin_134
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 46.837649402390866 0.25 47.087649402390866 ;
		END PORT
	END pin_134
	PIN pin_135
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 46.51792828685302 0.25 46.76792828685302 ;
		END PORT
	END pin_135
	PIN pin_136
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 46.198207171315175 0.25 46.448207171315175 ;
		END PORT
	END pin_136
	PIN pin_137
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 45.87848605577733 0.25 46.12848605577733 ;
		END PORT
	END pin_137
	PIN pin_138
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 45.558764940239485 0.25 45.808764940239485 ;
		END PORT
	END pin_138
	PIN pin_139
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 45.23904382470164 0.25 45.48904382470164 ;
		END PORT
	END pin_139
	PIN pin_140
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 44.919322709163794 0.25 45.169322709163794 ;
		END PORT
	END pin_140
	PIN pin_141
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 44.59960159362595 0.25 44.84960159362595 ;
		END PORT
	END pin_141
	PIN pin_142
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 44.2798804780881 0.25 44.5298804780881 ;
		END PORT
	END pin_142
	PIN pin_143
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 43.96015936255026 0.25 44.21015936255026 ;
		END PORT
	END pin_143
	PIN pin_144
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 43.64043824701241 0.25 43.89043824701241 ;
		END PORT
	END pin_144
	PIN pin_145
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 43.32071713147457 0.25 43.57071713147457 ;
		END PORT
	END pin_145
	PIN pin_146
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 43.00099601593672 0.25 43.25099601593672 ;
		END PORT
	END pin_146
	PIN pin_147
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 42.681274900398876 0.25 42.931274900398876 ;
		END PORT
	END pin_147
	PIN pin_148
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 42.36155378486103 0.25 42.61155378486103 ;
		END PORT
	END pin_148
	PIN pin_149
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 42.041832669323185 0.25 42.291832669323185 ;
		END PORT
	END pin_149
	PIN pin_150
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 41.72211155378534 0.25 41.97211155378534 ;
		END PORT
	END pin_150
	PIN pin_151
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 41.402390438247494 0.25 41.652390438247494 ;
		END PORT
	END pin_151
	PIN pin_152
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 41.08266932270965 0.25 41.33266932270965 ;
		END PORT
	END pin_152
	PIN pin_153
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 40.7629482071718 0.25 41.0129482071718 ;
		END PORT
	END pin_153
	PIN pin_154
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 40.44322709163396 0.25 40.69322709163396 ;
		END PORT
	END pin_154
	PIN pin_155
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 40.12350597609611 0.25 40.37350597609611 ;
		END PORT
	END pin_155
	PIN pin_156
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 39.80378486055827 0.25 40.05378486055827 ;
		END PORT
	END pin_156
	PIN pin_157
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 39.48406374502042 0.25 39.73406374502042 ;
		END PORT
	END pin_157
	PIN pin_158
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 39.164342629482576 0.25 39.414342629482576 ;
		END PORT
	END pin_158
	PIN pin_159
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 38.84462151394473 0.25 39.09462151394473 ;
		END PORT
	END pin_159
	PIN pin_160
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 38.524900398406885 0.25 38.774900398406885 ;
		END PORT
	END pin_160
	PIN pin_161
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 38.20517928286904 0.25 38.45517928286904 ;
		END PORT
	END pin_161
	PIN pin_162
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 37.885458167331194 0.25 38.135458167331194 ;
		END PORT
	END pin_162
	PIN pin_163
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 37.56573705179335 0.25 37.81573705179335 ;
		END PORT
	END pin_163
	PIN pin_164
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 37.2460159362555 0.25 37.4960159362555 ;
		END PORT
	END pin_164
	PIN pin_165
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 36.92629482071766 0.25 37.17629482071766 ;
		END PORT
	END pin_165
	PIN pin_166
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 36.60657370517981 0.25 36.85657370517981 ;
		END PORT
	END pin_166
	PIN pin_167
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 36.28685258964197 0.25 36.53685258964197 ;
		END PORT
	END pin_167
	PIN pin_168
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 35.96713147410412 0.25 36.21713147410412 ;
		END PORT
	END pin_168
	PIN pin_169
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 35.647410358566276 0.25 35.897410358566276 ;
		END PORT
	END pin_169
	PIN pin_170
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 35.32768924302843 0.25 35.57768924302843 ;
		END PORT
	END pin_170
	PIN pin_171
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 35.007968127490585 0.25 35.257968127490585 ;
		END PORT
	END pin_171
	PIN pin_172
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 34.68824701195274 0.25 34.93824701195274 ;
		END PORT
	END pin_172
	PIN pin_173
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 34.368525896414894 0.25 34.618525896414894 ;
		END PORT
	END pin_173
	PIN pin_174
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 34.04880478087705 0.25 34.29880478087705 ;
		END PORT
	END pin_174
	PIN pin_175
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 33.7290836653392 0.25 33.9790836653392 ;
		END PORT
	END pin_175
	PIN pin_176
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 33.40936254980136 0.25 33.65936254980136 ;
		END PORT
	END pin_176
	PIN pin_177
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 33.08964143426351 0.25 33.33964143426351 ;
		END PORT
	END pin_177
	PIN pin_178
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 32.76992031872567 0.25 33.01992031872567 ;
		END PORT
	END pin_178
	PIN pin_179
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 32.45019920318782 0.25 32.70019920318782 ;
		END PORT
	END pin_179
	PIN pin_180
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 32.130478087649976 0.25 32.380478087649976 ;
		END PORT
	END pin_180
	PIN pin_181
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 31.81075697211213 0.25 32.06075697211213 ;
		END PORT
	END pin_181
	PIN pin_182
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 31.491035856574282 0.25 31.741035856574282 ;
		END PORT
	END pin_182
	PIN pin_183
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 31.171314741036433 0.25 31.421314741036433 ;
		END PORT
	END pin_183
	PIN pin_184
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 30.851593625498584 0.25 31.101593625498584 ;
		END PORT
	END pin_184
	PIN pin_185
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 30.531872509960735 0.25 30.781872509960735 ;
		END PORT
	END pin_185
	PIN pin_186
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 30.212151394422886 0.25 30.462151394422886 ;
		END PORT
	END pin_186
	PIN pin_187
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 29.892430278885037 0.25 30.142430278885037 ;
		END PORT
	END pin_187
	PIN pin_188
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 29.572709163347188 0.25 29.822709163347188 ;
		END PORT
	END pin_188
	PIN pin_189
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 29.25298804780934 0.25 29.50298804780934 ;
		END PORT
	END pin_189
	PIN pin_190
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 28.93326693227149 0.25 29.18326693227149 ;
		END PORT
	END pin_190
	PIN pin_191
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 28.61354581673364 0.25 28.86354581673364 ;
		END PORT
	END pin_191
	PIN pin_192
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 28.293824701195792 0.25 28.543824701195792 ;
		END PORT
	END pin_192
	PIN pin_193
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 27.974103585657943 0.25 28.224103585657943 ;
		END PORT
	END pin_193
	PIN pin_194
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 27.654382470120094 0.25 27.904382470120094 ;
		END PORT
	END pin_194
	PIN pin_195
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 27.334661354582245 0.25 27.584661354582245 ;
		END PORT
	END pin_195
	PIN pin_196
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 27.014940239044396 0.25 27.264940239044396 ;
		END PORT
	END pin_196
	PIN pin_197
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 26.695219123506547 0.25 26.945219123506547 ;
		END PORT
	END pin_197
	PIN pin_198
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 26.375498007968698 0.25 26.625498007968698 ;
		END PORT
	END pin_198
	PIN pin_199
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 26.05577689243085 0.25 26.30577689243085 ;
		END PORT
	END pin_199
	PIN pin_200
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 25.736055776893 0.25 25.986055776893 ;
		END PORT
	END pin_200
	PIN pin_201
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 25.41633466135515 0.25 25.66633466135515 ;
		END PORT
	END pin_201
	PIN pin_202
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 25.096613545817302 0.25 25.346613545817302 ;
		END PORT
	END pin_202
	PIN pin_203
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 24.776892430279453 0.25 25.026892430279453 ;
		END PORT
	END pin_203
	PIN pin_204
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 24.457171314741604 0.25 24.707171314741604 ;
		END PORT
	END pin_204
	PIN pin_205
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 24.137450199203755 0.25 24.387450199203755 ;
		END PORT
	END pin_205
	PIN pin_206
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 23.817729083665906 0.25 24.067729083665906 ;
		END PORT
	END pin_206
	PIN pin_207
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 23.498007968128057 0.25 23.748007968128057 ;
		END PORT
	END pin_207
	PIN pin_208
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 23.178286852590208 0.25 23.428286852590208 ;
		END PORT
	END pin_208
	PIN pin_209
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 22.85856573705236 0.25 23.10856573705236 ;
		END PORT
	END pin_209
	PIN pin_210
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 22.53884462151451 0.25 22.78884462151451 ;
		END PORT
	END pin_210
	PIN pin_211
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 22.21912350597666 0.25 22.46912350597666 ;
		END PORT
	END pin_211
	PIN pin_212
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 21.899402390438812 0.25 22.149402390438812 ;
		END PORT
	END pin_212
	PIN pin_213
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 21.579681274900963 0.25 21.829681274900963 ;
		END PORT
	END pin_213
	PIN pin_214
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 21.259960159363114 0.25 21.509960159363114 ;
		END PORT
	END pin_214
	PIN pin_215
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 20.940239043825265 0.25 21.190239043825265 ;
		END PORT
	END pin_215
	PIN pin_216
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 20.620517928287416 0.25 20.870517928287416 ;
		END PORT
	END pin_216
	PIN pin_217
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 20.300796812749567 0.25 20.550796812749567 ;
		END PORT
	END pin_217
	PIN pin_218
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 19.98107569721172 0.25 20.23107569721172 ;
		END PORT
	END pin_218
	PIN pin_219
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 19.66135458167387 0.25 19.91135458167387 ;
		END PORT
	END pin_219
	PIN pin_220
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 19.34163346613602 0.25 19.59163346613602 ;
		END PORT
	END pin_220
	PIN pin_221
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 19.02191235059817 0.25 19.27191235059817 ;
		END PORT
	END pin_221
	PIN pin_222
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 18.702191235060322 0.25 18.952191235060322 ;
		END PORT
	END pin_222
	PIN pin_223
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 18.382470119522473 0.25 18.632470119522473 ;
		END PORT
	END pin_223
	PIN pin_224
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 18.062749003984624 0.25 18.312749003984624 ;
		END PORT
	END pin_224
	PIN pin_225
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 17.743027888446775 0.25 17.993027888446775 ;
		END PORT
	END pin_225
	PIN pin_226
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 17.423306772908926 0.25 17.673306772908926 ;
		END PORT
	END pin_226
	PIN pin_227
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 17.103585657371077 0.25 17.353585657371077 ;
		END PORT
	END pin_227
	PIN pin_228
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 16.78386454183323 0.25 17.03386454183323 ;
		END PORT
	END pin_228
	PIN pin_229
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 16.46414342629538 0.25 16.71414342629538 ;
		END PORT
	END pin_229
	PIN pin_230
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 16.14442231075753 0.25 16.39442231075753 ;
		END PORT
	END pin_230
	PIN pin_231
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 15.824701195219681 0.25 16.07470119521968 ;
		END PORT
	END pin_231
	PIN pin_232
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 15.504980079681832 0.25 15.754980079681832 ;
		END PORT
	END pin_232
	PIN pin_233
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 15.185258964143983 0.25 15.435258964143983 ;
		END PORT
	END pin_233
	PIN pin_234
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 14.865537848606134 0.25 15.115537848606134 ;
		END PORT
	END pin_234
	PIN pin_235
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 14.545816733068285 0.25 14.795816733068285 ;
		END PORT
	END pin_235
	PIN pin_236
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 14.226095617530436 0.25 14.476095617530436 ;
		END PORT
	END pin_236
	PIN pin_237
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 13.906374501992588 0.25 14.156374501992588 ;
		END PORT
	END pin_237
	PIN pin_238
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 13.586653386454739 0.25 13.836653386454739 ;
		END PORT
	END pin_238
	PIN pin_239
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 13.26693227091689 0.25 13.51693227091689 ;
		END PORT
	END pin_239
	PIN pin_240
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 12.94721115537904 0.25 13.19721115537904 ;
		END PORT
	END pin_240
	PIN pin_241
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 12.627490039841192 0.25 12.877490039841192 ;
		END PORT
	END pin_241
	PIN pin_242
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 12.307768924303343 0.25 12.557768924303343 ;
		END PORT
	END pin_242
	PIN pin_243
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 11.988047808765494 0.25 12.238047808765494 ;
		END PORT
	END pin_243
	PIN pin_244
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 11.668326693227645 0.25 11.918326693227645 ;
		END PORT
	END pin_244
	PIN pin_245
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 11.348605577689796 0.25 11.598605577689796 ;
		END PORT
	END pin_245
	PIN pin_246
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 11.028884462151947 0.25 11.278884462151947 ;
		END PORT
	END pin_246
	PIN pin_247
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 10.709163346614098 0.25 10.959163346614098 ;
		END PORT
	END pin_247
	PIN pin_248
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 10.389442231076249 0.25 10.639442231076249 ;
		END PORT
	END pin_248
	PIN pin_249
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 10.0697211155384 0.25 10.3197211155384 ;
		END PORT
	END pin_249
	PIN pin_250
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.069721115537849 100 10.319721115537849 ;
		END PORT
	END pin_250
	PIN pin_251
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.389442231075698 100 10.639442231075698 ;
		END PORT
	END pin_251
	PIN pin_252
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.709163346613547 100 10.959163346613547 ;
		END PORT
	END pin_252
	PIN pin_253
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.028884462151396 100 11.278884462151396 ;
		END PORT
	END pin_253
	PIN pin_254
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.348605577689245 100 11.598605577689245 ;
		END PORT
	END pin_254
	PIN pin_255
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.668326693227094 100 11.918326693227094 ;
		END PORT
	END pin_255
	PIN pin_256
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.988047808764943 100 12.238047808764943 ;
		END PORT
	END pin_256
	PIN pin_257
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.307768924302792 100 12.557768924302792 ;
		END PORT
	END pin_257
	PIN pin_258
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.627490039840641 100 12.877490039840641 ;
		END PORT
	END pin_258
	PIN pin_259
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.94721115537849 100 13.19721115537849 ;
		END PORT
	END pin_259
	PIN pin_260
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.266932270916339 100 13.516932270916339 ;
		END PORT
	END pin_260
	PIN pin_261
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.586653386454188 100 13.836653386454188 ;
		END PORT
	END pin_261
	PIN pin_262
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.906374501992037 100 14.156374501992037 ;
		END PORT
	END pin_262
	PIN pin_263
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.226095617529886 100 14.476095617529886 ;
		END PORT
	END pin_263
	PIN pin_264
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.545816733067735 100 14.795816733067735 ;
		END PORT
	END pin_264
	PIN pin_265
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.865537848605584 100 15.115537848605584 ;
		END PORT
	END pin_265
	PIN pin_266
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.185258964143433 100 15.435258964143433 ;
		END PORT
	END pin_266
	PIN pin_267
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.504980079681282 100 15.754980079681282 ;
		END PORT
	END pin_267
	PIN pin_268
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.82470119521913 100 16.07470119521913 ;
		END PORT
	END pin_268
	PIN pin_269
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.14442231075698 100 16.39442231075698 ;
		END PORT
	END pin_269
	PIN pin_270
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.46414342629483 100 16.71414342629483 ;
		END PORT
	END pin_270
	PIN pin_271
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.783864541832678 100 17.033864541832678 ;
		END PORT
	END pin_271
	PIN pin_272
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.103585657370527 100 17.353585657370527 ;
		END PORT
	END pin_272
	PIN pin_273
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.423306772908376 100 17.673306772908376 ;
		END PORT
	END pin_273
	PIN pin_274
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.743027888446225 100 17.993027888446225 ;
		END PORT
	END pin_274
	PIN pin_275
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.062749003984074 100 18.312749003984074 ;
		END PORT
	END pin_275
	PIN pin_276
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.382470119521923 100 18.632470119521923 ;
		END PORT
	END pin_276
	PIN pin_277
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.70219123505977 100 18.95219123505977 ;
		END PORT
	END pin_277
	PIN pin_278
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.02191235059762 100 19.27191235059762 ;
		END PORT
	END pin_278
	PIN pin_279
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.34163346613547 100 19.59163346613547 ;
		END PORT
	END pin_279
	PIN pin_280
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.66135458167332 100 19.91135458167332 ;
		END PORT
	END pin_280
	PIN pin_281
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.981075697211168 100 20.231075697211168 ;
		END PORT
	END pin_281
	PIN pin_282
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.300796812749017 100 20.550796812749017 ;
		END PORT
	END pin_282
	PIN pin_283
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.620517928286866 100 20.870517928286866 ;
		END PORT
	END pin_283
	PIN pin_284
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.940239043824715 100 21.190239043824715 ;
		END PORT
	END pin_284
	PIN pin_285
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.259960159362564 100 21.509960159362564 ;
		END PORT
	END pin_285
	PIN pin_286
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.579681274900413 100 21.829681274900413 ;
		END PORT
	END pin_286
	PIN pin_287
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.89940239043826 100 22.14940239043826 ;
		END PORT
	END pin_287
	PIN pin_288
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.21912350597611 100 22.46912350597611 ;
		END PORT
	END pin_288
	PIN pin_289
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.53884462151396 100 22.78884462151396 ;
		END PORT
	END pin_289
	PIN pin_290
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.85856573705181 100 23.10856573705181 ;
		END PORT
	END pin_290
	PIN pin_291
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.178286852589657 100 23.428286852589657 ;
		END PORT
	END pin_291
	PIN pin_292
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.498007968127506 100 23.748007968127506 ;
		END PORT
	END pin_292
	PIN pin_293
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.817729083665355 100 24.067729083665355 ;
		END PORT
	END pin_293
	PIN pin_294
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.137450199203204 100 24.387450199203204 ;
		END PORT
	END pin_294
	PIN pin_295
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.457171314741053 100 24.707171314741053 ;
		END PORT
	END pin_295
	PIN pin_296
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.776892430278902 100 25.026892430278902 ;
		END PORT
	END pin_296
	PIN pin_297
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.09661354581675 100 25.34661354581675 ;
		END PORT
	END pin_297
	PIN pin_298
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.4163346613546 100 25.6663346613546 ;
		END PORT
	END pin_298
	PIN pin_299
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.73605577689245 100 25.98605577689245 ;
		END PORT
	END pin_299
	PIN pin_300
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.0557768924303 100 26.3057768924303 ;
		END PORT
	END pin_300
	PIN pin_301
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.375498007968147 100 26.625498007968147 ;
		END PORT
	END pin_301
	PIN pin_302
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.695219123505996 100 26.945219123505996 ;
		END PORT
	END pin_302
	PIN pin_303
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.014940239043845 100 27.264940239043845 ;
		END PORT
	END pin_303
	PIN pin_304
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.334661354581694 100 27.584661354581694 ;
		END PORT
	END pin_304
	PIN pin_305
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.654382470119543 100 27.904382470119543 ;
		END PORT
	END pin_305
	PIN pin_306
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.974103585657392 100 28.224103585657392 ;
		END PORT
	END pin_306
	PIN pin_307
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.29382470119524 100 28.54382470119524 ;
		END PORT
	END pin_307
	PIN pin_308
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.61354581673309 100 28.86354581673309 ;
		END PORT
	END pin_308
	PIN pin_309
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.93326693227094 100 29.18326693227094 ;
		END PORT
	END pin_309
	PIN pin_310
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.25298804780879 100 29.50298804780879 ;
		END PORT
	END pin_310
	PIN pin_311
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.572709163346637 100 29.822709163346637 ;
		END PORT
	END pin_311
	PIN pin_312
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.892430278884486 100 30.142430278884486 ;
		END PORT
	END pin_312
	PIN pin_313
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.212151394422335 100 30.462151394422335 ;
		END PORT
	END pin_313
	PIN pin_314
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.531872509960184 100 30.781872509960184 ;
		END PORT
	END pin_314
	PIN pin_315
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.851593625498033 100 31.101593625498033 ;
		END PORT
	END pin_315
	PIN pin_316
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.171314741035882 100 31.421314741035882 ;
		END PORT
	END pin_316
	PIN pin_317
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.49103585657373 100 31.74103585657373 ;
		END PORT
	END pin_317
	PIN pin_318
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.81075697211158 100 32.06075697211158 ;
		END PORT
	END pin_318
	PIN pin_319
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.13047808764942 100 32.38047808764942 ;
		END PORT
	END pin_319
	PIN pin_320
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.45019920318727 100 32.70019920318727 ;
		END PORT
	END pin_320
	PIN pin_321
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.76992031872511 100 33.01992031872511 ;
		END PORT
	END pin_321
	PIN pin_322
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.08964143426296 100 33.33964143426296 ;
		END PORT
	END pin_322
	PIN pin_323
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.409362549800804 100 33.659362549800804 ;
		END PORT
	END pin_323
	PIN pin_324
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.72908366533865 100 33.97908366533865 ;
		END PORT
	END pin_324
	PIN pin_325
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.048804780876495 100 34.298804780876495 ;
		END PORT
	END pin_325
	PIN pin_326
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.36852589641434 100 34.61852589641434 ;
		END PORT
	END pin_326
	PIN pin_327
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.688247011952186 100 34.938247011952186 ;
		END PORT
	END pin_327
	PIN pin_328
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.00796812749003 100 35.25796812749003 ;
		END PORT
	END pin_328
	PIN pin_329
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.327689243027876 100 35.577689243027876 ;
		END PORT
	END pin_329
	PIN pin_330
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.64741035856572 100 35.89741035856572 ;
		END PORT
	END pin_330
	PIN pin_331
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.96713147410357 100 36.21713147410357 ;
		END PORT
	END pin_331
	PIN pin_332
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.28685258964141 100 36.53685258964141 ;
		END PORT
	END pin_332
	PIN pin_333
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.60657370517926 100 36.85657370517926 ;
		END PORT
	END pin_333
	PIN pin_334
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.926294820717104 100 37.176294820717104 ;
		END PORT
	END pin_334
	PIN pin_335
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.24601593625495 100 37.49601593625495 ;
		END PORT
	END pin_335
	PIN pin_336
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.565737051792794 100 37.815737051792794 ;
		END PORT
	END pin_336
	PIN pin_337
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.88545816733064 100 38.13545816733064 ;
		END PORT
	END pin_337
	PIN pin_338
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.205179282868485 100 38.455179282868485 ;
		END PORT
	END pin_338
	PIN pin_339
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.52490039840633 100 38.77490039840633 ;
		END PORT
	END pin_339
	PIN pin_340
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.844621513944176 100 39.094621513944176 ;
		END PORT
	END pin_340
	PIN pin_341
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.16434262948202 100 39.41434262948202 ;
		END PORT
	END pin_341
	PIN pin_342
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.48406374501987 100 39.73406374501987 ;
		END PORT
	END pin_342
	PIN pin_343
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.80378486055771 100 40.05378486055771 ;
		END PORT
	END pin_343
	PIN pin_344
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.12350597609556 100 40.37350597609556 ;
		END PORT
	END pin_344
	PIN pin_345
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.4432270916334 100 40.6932270916334 ;
		END PORT
	END pin_345
	PIN pin_346
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.76294820717125 100 41.01294820717125 ;
		END PORT
	END pin_346
	PIN pin_347
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.082669322709094 100 41.332669322709094 ;
		END PORT
	END pin_347
	PIN pin_348
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.40239043824694 100 41.65239043824694 ;
		END PORT
	END pin_348
	PIN pin_349
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.722111553784785 100 41.972111553784785 ;
		END PORT
	END pin_349
	PIN pin_350
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.04183266932263 100 42.29183266932263 ;
		END PORT
	END pin_350
	PIN pin_351
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.361553784860476 100 42.611553784860476 ;
		END PORT
	END pin_351
	PIN pin_352
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.68127490039832 100 42.93127490039832 ;
		END PORT
	END pin_352
	PIN pin_353
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.00099601593617 100 43.25099601593617 ;
		END PORT
	END pin_353
	PIN pin_354
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.32071713147401 100 43.57071713147401 ;
		END PORT
	END pin_354
	PIN pin_355
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.64043824701186 100 43.89043824701186 ;
		END PORT
	END pin_355
	PIN pin_356
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.9601593625497 100 44.2101593625497 ;
		END PORT
	END pin_356
	PIN pin_357
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.27988047808755 100 44.52988047808755 ;
		END PORT
	END pin_357
	PIN pin_358
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.599601593625394 100 44.849601593625394 ;
		END PORT
	END pin_358
	PIN pin_359
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.91932270916324 100 45.16932270916324 ;
		END PORT
	END pin_359
	PIN pin_360
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.239043824701085 100 45.489043824701085 ;
		END PORT
	END pin_360
	PIN pin_361
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.55876494023893 100 45.80876494023893 ;
		END PORT
	END pin_361
	PIN pin_362
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.878486055776776 100 46.128486055776776 ;
		END PORT
	END pin_362
	PIN pin_363
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.19820717131462 100 46.44820717131462 ;
		END PORT
	END pin_363
	PIN pin_364
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.51792828685247 100 46.76792828685247 ;
		END PORT
	END pin_364
	PIN pin_365
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.83764940239031 100 47.08764940239031 ;
		END PORT
	END pin_365
	PIN pin_366
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.15737051792816 100 47.40737051792816 ;
		END PORT
	END pin_366
	PIN pin_367
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.477091633466 100 47.727091633466 ;
		END PORT
	END pin_367
	PIN pin_368
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.79681274900385 100 48.04681274900385 ;
		END PORT
	END pin_368
	PIN pin_369
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.116533864541694 100 48.366533864541694 ;
		END PORT
	END pin_369
	PIN pin_370
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.43625498007954 100 48.68625498007954 ;
		END PORT
	END pin_370
	PIN pin_371
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.755976095617385 100 49.005976095617385 ;
		END PORT
	END pin_371
	PIN pin_372
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.07569721115523 100 49.32569721115523 ;
		END PORT
	END pin_372
	PIN pin_373
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.395418326693076 100 49.645418326693076 ;
		END PORT
	END pin_373
	PIN pin_374
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.71513944223092 100 49.96513944223092 ;
		END PORT
	END pin_374
	PIN pin_375
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.034860557768766 100 50.284860557768766 ;
		END PORT
	END pin_375
	PIN pin_376
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.35458167330661 100 50.60458167330661 ;
		END PORT
	END pin_376
	PIN pin_377
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.67430278884446 100 50.92430278884446 ;
		END PORT
	END pin_377
	PIN pin_378
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.9940239043823 100 51.2440239043823 ;
		END PORT
	END pin_378
	PIN pin_379
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.31374501992015 100 51.56374501992015 ;
		END PORT
	END pin_379
	PIN pin_380
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.633466135457994 100 51.883466135457994 ;
		END PORT
	END pin_380
	PIN pin_381
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.95318725099584 100 52.20318725099584 ;
		END PORT
	END pin_381
	PIN pin_382
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.272908366533684 100 52.522908366533684 ;
		END PORT
	END pin_382
	PIN pin_383
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.59262948207153 100 52.84262948207153 ;
		END PORT
	END pin_383
	PIN pin_384
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.912350597609375 100 53.162350597609375 ;
		END PORT
	END pin_384
	PIN pin_385
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.23207171314722 100 53.48207171314722 ;
		END PORT
	END pin_385
	PIN pin_386
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.551792828685066 100 53.801792828685066 ;
		END PORT
	END pin_386
	PIN pin_387
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.87151394422291 100 54.12151394422291 ;
		END PORT
	END pin_387
	PIN pin_388
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.19123505976076 100 54.44123505976076 ;
		END PORT
	END pin_388
	PIN pin_389
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.5109561752986 100 54.7609561752986 ;
		END PORT
	END pin_389
	PIN pin_390
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.83067729083645 100 55.08067729083645 ;
		END PORT
	END pin_390
	PIN pin_391
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.15039840637429 100 55.40039840637429 ;
		END PORT
	END pin_391
	PIN pin_392
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.47011952191214 100 55.72011952191214 ;
		END PORT
	END pin_392
	PIN pin_393
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.789840637449984 100 56.039840637449984 ;
		END PORT
	END pin_393
	PIN pin_394
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.10956175298783 100 56.35956175298783 ;
		END PORT
	END pin_394
	PIN pin_395
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.429282868525675 100 56.679282868525675 ;
		END PORT
	END pin_395
	PIN pin_396
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.74900398406352 100 56.99900398406352 ;
		END PORT
	END pin_396
	PIN pin_397
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.068725099601366 100 57.318725099601366 ;
		END PORT
	END pin_397
	PIN pin_398
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.38844621513921 100 57.63844621513921 ;
		END PORT
	END pin_398
	PIN pin_399
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.70816733067706 100 57.95816733067706 ;
		END PORT
	END pin_399
	PIN pin_400
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.0278884462149 100 58.2778884462149 ;
		END PORT
	END pin_400
	PIN pin_401
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.34760956175275 100 58.59760956175275 ;
		END PORT
	END pin_401
	PIN pin_402
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.66733067729059 100 58.91733067729059 ;
		END PORT
	END pin_402
	PIN pin_403
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.98705179282844 100 59.23705179282844 ;
		END PORT
	END pin_403
	PIN pin_404
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.306772908366284 100 59.556772908366284 ;
		END PORT
	END pin_404
	PIN pin_405
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.62649402390413 100 59.87649402390413 ;
		END PORT
	END pin_405
	PIN pin_406
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.946215139441975 100 60.196215139441975 ;
		END PORT
	END pin_406
	PIN pin_407
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.26593625497982 100 60.51593625497982 ;
		END PORT
	END pin_407
	PIN pin_408
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.585657370517666 100 60.835657370517666 ;
		END PORT
	END pin_408
	PIN pin_409
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.90537848605551 100 61.15537848605551 ;
		END PORT
	END pin_409
	PIN pin_410
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.22509960159336 100 61.47509960159336 ;
		END PORT
	END pin_410
	PIN pin_411
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.5448207171312 100 61.7948207171312 ;
		END PORT
	END pin_411
	PIN pin_412
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.86454183266905 100 62.11454183266905 ;
		END PORT
	END pin_412
	PIN pin_413
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.18426294820689 100 62.43426294820689 ;
		END PORT
	END pin_413
	PIN pin_414
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.50398406374474 100 62.75398406374474 ;
		END PORT
	END pin_414
	PIN pin_415
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.823705179282584 100 63.073705179282584 ;
		END PORT
	END pin_415
	PIN pin_416
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.14342629482043 100 63.39342629482043 ;
		END PORT
	END pin_416
	PIN pin_417
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.463147410358275 100 63.713147410358275 ;
		END PORT
	END pin_417
	PIN pin_418
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.78286852589612 100 64.03286852589612 ;
		END PORT
	END pin_418
	PIN pin_419
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.10258964143397 100 64.35258964143397 ;
		END PORT
	END pin_419
	PIN pin_420
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.42231075697181 100 64.67231075697181 ;
		END PORT
	END pin_420
	PIN pin_421
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.74203187250966 100 64.99203187250966 ;
		END PORT
	END pin_421
	PIN pin_422
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.0617529880475 100 65.3117529880475 ;
		END PORT
	END pin_422
	PIN pin_423
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.38147410358535 100 65.63147410358535 ;
		END PORT
	END pin_423
	PIN pin_424
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.70119521912319 100 65.95119521912319 ;
		END PORT
	END pin_424
	PIN pin_425
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.02091633466104 100 66.27091633466104 ;
		END PORT
	END pin_425
	PIN pin_426
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.34063745019888 100 66.59063745019888 ;
		END PORT
	END pin_426
	PIN pin_427
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.66035856573673 100 66.91035856573673 ;
		END PORT
	END pin_427
	PIN pin_428
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.98007968127457 100 67.23007968127457 ;
		END PORT
	END pin_428
	PIN pin_429
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.29980079681242 100 67.54980079681242 ;
		END PORT
	END pin_429
	PIN pin_430
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.61952191235027 100 67.86952191235027 ;
		END PORT
	END pin_430
	PIN pin_431
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.93924302788811 100 68.18924302788811 ;
		END PORT
	END pin_431
	PIN pin_432
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.25896414342596 100 68.50896414342596 ;
		END PORT
	END pin_432
	PIN pin_433
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.5786852589638 100 68.8286852589638 ;
		END PORT
	END pin_433
	PIN pin_434
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.89840637450165 100 69.14840637450165 ;
		END PORT
	END pin_434
	PIN pin_435
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.21812749003949 100 69.46812749003949 ;
		END PORT
	END pin_435
	PIN pin_436
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.53784860557734 100 69.78784860557734 ;
		END PORT
	END pin_436
	PIN pin_437
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.85756972111518 100 70.10756972111518 ;
		END PORT
	END pin_437
	PIN pin_438
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.17729083665303 100 70.42729083665303 ;
		END PORT
	END pin_438
	PIN pin_439
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.49701195219087 100 70.74701195219087 ;
		END PORT
	END pin_439
	PIN pin_440
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.81673306772872 100 71.06673306772872 ;
		END PORT
	END pin_440
	PIN pin_441
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.13645418326657 100 71.38645418326657 ;
		END PORT
	END pin_441
	PIN pin_442
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.45617529880441 100 71.70617529880441 ;
		END PORT
	END pin_442
	PIN pin_443
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.77589641434226 100 72.02589641434226 ;
		END PORT
	END pin_443
	PIN pin_444
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.0956175298801 100 72.3456175298801 ;
		END PORT
	END pin_444
	PIN pin_445
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.41533864541795 100 72.66533864541795 ;
		END PORT
	END pin_445
	PIN pin_446
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.73505976095579 100 72.98505976095579 ;
		END PORT
	END pin_446
	PIN pin_447
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.05478087649364 100 73.30478087649364 ;
		END PORT
	END pin_447
	PIN pin_448
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.37450199203148 100 73.62450199203148 ;
		END PORT
	END pin_448
	PIN pin_449
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.69422310756933 100 73.94422310756933 ;
		END PORT
	END pin_449
	PIN pin_450
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.01394422310717 100 74.26394422310717 ;
		END PORT
	END pin_450
	PIN pin_451
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.33366533864502 100 74.58366533864502 ;
		END PORT
	END pin_451
	PIN pin_452
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.65338645418286 100 74.90338645418286 ;
		END PORT
	END pin_452
	PIN pin_453
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.97310756972071 100 75.22310756972071 ;
		END PORT
	END pin_453
	PIN pin_454
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.29282868525856 100 75.54282868525856 ;
		END PORT
	END pin_454
	PIN pin_455
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.6125498007964 100 75.8625498007964 ;
		END PORT
	END pin_455
	PIN pin_456
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.93227091633425 100 76.18227091633425 ;
		END PORT
	END pin_456
	PIN pin_457
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.25199203187209 100 76.50199203187209 ;
		END PORT
	END pin_457
	PIN pin_458
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.57171314740994 100 76.82171314740994 ;
		END PORT
	END pin_458
	PIN pin_459
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.89143426294778 100 77.14143426294778 ;
		END PORT
	END pin_459
	PIN pin_460
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.21115537848563 100 77.46115537848563 ;
		END PORT
	END pin_460
	PIN pin_461
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.53087649402347 100 77.78087649402347 ;
		END PORT
	END pin_461
	PIN pin_462
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.85059760956132 100 78.10059760956132 ;
		END PORT
	END pin_462
	PIN pin_463
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.17031872509916 100 78.42031872509916 ;
		END PORT
	END pin_463
	PIN pin_464
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.49003984063701 100 78.74003984063701 ;
		END PORT
	END pin_464
	PIN pin_465
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.80976095617486 100 79.05976095617486 ;
		END PORT
	END pin_465
	PIN pin_466
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.1294820717127 100 79.3794820717127 ;
		END PORT
	END pin_466
	PIN pin_467
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.44920318725055 100 79.69920318725055 ;
		END PORT
	END pin_467
	PIN pin_468
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.76892430278839 100 80.01892430278839 ;
		END PORT
	END pin_468
	PIN pin_469
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.08864541832624 100 80.33864541832624 ;
		END PORT
	END pin_469
	PIN pin_470
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.40836653386408 100 80.65836653386408 ;
		END PORT
	END pin_470
	PIN pin_471
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.72808764940193 100 80.97808764940193 ;
		END PORT
	END pin_471
	PIN pin_472
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.04780876493977 100 81.29780876493977 ;
		END PORT
	END pin_472
	PIN pin_473
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.36752988047762 100 81.61752988047762 ;
		END PORT
	END pin_473
	PIN pin_474
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.68725099601546 100 81.93725099601546 ;
		END PORT
	END pin_474
	PIN pin_475
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.00697211155331 100 82.25697211155331 ;
		END PORT
	END pin_475
	PIN pin_476
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.32669322709116 100 82.57669322709116 ;
		END PORT
	END pin_476
	PIN pin_477
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.646414342629 100 82.896414342629 ;
		END PORT
	END pin_477
	PIN pin_478
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.96613545816685 100 83.21613545816685 ;
		END PORT
	END pin_478
	PIN pin_479
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.28585657370469 100 83.53585657370469 ;
		END PORT
	END pin_479
	PIN pin_480
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.60557768924254 100 83.85557768924254 ;
		END PORT
	END pin_480
	PIN pin_481
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.92529880478038 100 84.17529880478038 ;
		END PORT
	END pin_481
	PIN pin_482
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.24501992031823 100 84.49501992031823 ;
		END PORT
	END pin_482
	PIN pin_483
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.56474103585607 100 84.81474103585607 ;
		END PORT
	END pin_483
	PIN pin_484
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.88446215139392 100 85.13446215139392 ;
		END PORT
	END pin_484
	PIN pin_485
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.20418326693176 100 85.45418326693176 ;
		END PORT
	END pin_485
	PIN pin_486
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.52390438246961 100 85.77390438246961 ;
		END PORT
	END pin_486
	PIN pin_487
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.84362549800746 100 86.09362549800746 ;
		END PORT
	END pin_487
	PIN pin_488
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.1633466135453 100 86.4133466135453 ;
		END PORT
	END pin_488
	PIN pin_489
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.48306772908315 100 86.73306772908315 ;
		END PORT
	END pin_489
	PIN pin_490
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.80278884462099 100 87.05278884462099 ;
		END PORT
	END pin_490
	PIN pin_491
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.12250996015884 100 87.37250996015884 ;
		END PORT
	END pin_491
	PIN pin_492
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.44223107569668 100 87.69223107569668 ;
		END PORT
	END pin_492
	PIN pin_493
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.76195219123453 100 88.01195219123453 ;
		END PORT
	END pin_493
	PIN pin_494
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.08167330677237 100 88.33167330677237 ;
		END PORT
	END pin_494
	PIN pin_495
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.40139442231022 100 88.65139442231022 ;
		END PORT
	END pin_495
	PIN pin_496
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.72111553784806 100 88.97111553784806 ;
		END PORT
	END pin_496
	PIN pin_497
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.04083665338591 100 89.29083665338591 ;
		END PORT
	END pin_497
	PIN pin_498
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.36055776892375 100 89.61055776892375 ;
		END PORT
	END pin_498
	PIN pin_499
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.6802788844616 100 89.9302788844616 ;
		END PORT
	END pin_499
	PIN pin_500
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 89.68027888446215 99.75 89.93027888446215 100 ;
		END PORT
	END pin_500
	PIN pin_501
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.36055776892431 99.75 89.61055776892431 100 ;
		END PORT
	END pin_501
	PIN pin_502
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 89.04083665338646 99.75 89.29083665338646 100 ;
		END PORT
	END pin_502
	PIN pin_503
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.72111553784862 99.75 88.97111553784862 100 ;
		END PORT
	END pin_503
	PIN pin_504
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 88.40139442231077 99.75 88.65139442231077 100 ;
		END PORT
	END pin_504
	PIN pin_505
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.08167330677293 99.75 88.33167330677293 100 ;
		END PORT
	END pin_505
	PIN pin_506
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.76195219123508 99.75 88.01195219123508 100 ;
		END PORT
	END pin_506
	PIN pin_507
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 87.44223107569724 99.75 87.69223107569724 100 ;
		END PORT
	END pin_507
	PIN pin_508
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 87.12250996015939 99.75 87.37250996015939 100 ;
		END PORT
	END pin_508
	PIN pin_509
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.80278884462155 99.75 87.05278884462155 100 ;
		END PORT
	END pin_509
	PIN pin_510
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 86.4830677290837 99.75 86.7330677290837 100 ;
		END PORT
	END pin_510
	PIN pin_511
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 86.16334661354585 99.75 86.41334661354585 100 ;
		END PORT
	END pin_511
	PIN pin_512
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.84362549800801 99.75 86.09362549800801 100 ;
		END PORT
	END pin_512
	PIN pin_513
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 85.52390438247016 99.75 85.77390438247016 100 ;
		END PORT
	END pin_513
	PIN pin_514
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 85.20418326693232 99.75 85.45418326693232 100 ;
		END PORT
	END pin_514
	PIN pin_515
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 84.88446215139447 99.75 85.13446215139447 100 ;
		END PORT
	END pin_515
	PIN pin_516
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 84.56474103585663 99.75 84.81474103585663 100 ;
		END PORT
	END pin_516
	PIN pin_517
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 84.24501992031878 99.75 84.49501992031878 100 ;
		END PORT
	END pin_517
	PIN pin_518
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.92529880478094 99.75 84.17529880478094 100 ;
		END PORT
	END pin_518
	PIN pin_519
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 83.60557768924309 99.75 83.85557768924309 100 ;
		END PORT
	END pin_519
	PIN pin_520
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.28585657370525 99.75 83.53585657370525 100 ;
		END PORT
	END pin_520
	PIN pin_521
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.9661354581674 99.75 83.2161354581674 100 ;
		END PORT
	END pin_521
	PIN pin_522
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.64641434262955 99.75 82.89641434262955 100 ;
		END PORT
	END pin_522
	PIN pin_523
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.32669322709171 99.75 82.57669322709171 100 ;
		END PORT
	END pin_523
	PIN pin_524
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.00697211155386 99.75 82.25697211155386 100 ;
		END PORT
	END pin_524
	PIN pin_525
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.68725099601602 99.75 81.93725099601602 100 ;
		END PORT
	END pin_525
	PIN pin_526
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 81.36752988047817 99.75 81.61752988047817 100 ;
		END PORT
	END pin_526
	PIN pin_527
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.04780876494033 99.75 81.29780876494033 100 ;
		END PORT
	END pin_527
	PIN pin_528
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 80.72808764940248 99.75 80.97808764940248 100 ;
		END PORT
	END pin_528
	PIN pin_529
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 80.40836653386464 99.75 80.65836653386464 100 ;
		END PORT
	END pin_529
	PIN pin_530
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 80.08864541832679 99.75 80.33864541832679 100 ;
		END PORT
	END pin_530
	PIN pin_531
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.76892430278895 99.75 80.01892430278895 100 ;
		END PORT
	END pin_531
	PIN pin_532
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.4492031872511 99.75 79.6992031872511 100 ;
		END PORT
	END pin_532
	PIN pin_533
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.12948207171326 99.75 79.37948207171326 100 ;
		END PORT
	END pin_533
	PIN pin_534
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 78.80976095617541 99.75 79.05976095617541 100 ;
		END PORT
	END pin_534
	PIN pin_535
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 78.49003984063756 99.75 78.74003984063756 100 ;
		END PORT
	END pin_535
	PIN pin_536
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 78.17031872509972 99.75 78.42031872509972 100 ;
		END PORT
	END pin_536
	PIN pin_537
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.85059760956187 99.75 78.10059760956187 100 ;
		END PORT
	END pin_537
	PIN pin_538
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.53087649402403 99.75 77.78087649402403 100 ;
		END PORT
	END pin_538
	PIN pin_539
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 77.21115537848618 99.75 77.46115537848618 100 ;
		END PORT
	END pin_539
	PIN pin_540
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.89143426294834 99.75 77.14143426294834 100 ;
		END PORT
	END pin_540
	PIN pin_541
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 76.57171314741049 99.75 76.82171314741049 100 ;
		END PORT
	END pin_541
	PIN pin_542
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 76.25199203187265 99.75 76.50199203187265 100 ;
		END PORT
	END pin_542
	PIN pin_543
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 75.9322709163348 99.75 76.1822709163348 100 ;
		END PORT
	END pin_543
	PIN pin_544
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.61254980079696 99.75 75.86254980079696 100 ;
		END PORT
	END pin_544
	PIN pin_545
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 75.29282868525911 99.75 75.54282868525911 100 ;
		END PORT
	END pin_545
	PIN pin_546
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.97310756972126 99.75 75.22310756972126 100 ;
		END PORT
	END pin_546
	PIN pin_547
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 74.65338645418342 99.75 74.90338645418342 100 ;
		END PORT
	END pin_547
	PIN pin_548
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 74.33366533864557 99.75 74.58366533864557 100 ;
		END PORT
	END pin_548
	PIN pin_549
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.01394422310773 99.75 74.26394422310773 100 ;
		END PORT
	END pin_549
	PIN pin_550
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.69422310756988 99.75 73.94422310756988 100 ;
		END PORT
	END pin_550
	PIN pin_551
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.37450199203204 99.75 73.62450199203204 100 ;
		END PORT
	END pin_551
	PIN pin_552
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 73.05478087649419 99.75 73.30478087649419 100 ;
		END PORT
	END pin_552
	PIN pin_553
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 72.73505976095635 99.75 72.98505976095635 100 ;
		END PORT
	END pin_553
	PIN pin_554
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 72.4153386454185 99.75 72.6653386454185 100 ;
		END PORT
	END pin_554
	PIN pin_555
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 72.09561752988066 99.75 72.34561752988066 100 ;
		END PORT
	END pin_555
	PIN pin_556
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 71.77589641434281 99.75 72.02589641434281 100 ;
		END PORT
	END pin_556
	PIN pin_557
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 71.45617529880496 99.75 71.70617529880496 100 ;
		END PORT
	END pin_557
	PIN pin_558
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 71.13645418326712 99.75 71.38645418326712 100 ;
		END PORT
	END pin_558
	PIN pin_559
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 70.81673306772927 99.75 71.06673306772927 100 ;
		END PORT
	END pin_559
	PIN pin_560
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 70.49701195219143 99.75 70.74701195219143 100 ;
		END PORT
	END pin_560
	PIN pin_561
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 70.17729083665358 99.75 70.42729083665358 100 ;
		END PORT
	END pin_561
	PIN pin_562
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 69.85756972111574 99.75 70.10756972111574 100 ;
		END PORT
	END pin_562
	PIN pin_563
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 69.53784860557789 99.75 69.78784860557789 100 ;
		END PORT
	END pin_563
	PIN pin_564
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 69.21812749004005 99.75 69.46812749004005 100 ;
		END PORT
	END pin_564
	PIN pin_565
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.8984063745022 99.75 69.1484063745022 100 ;
		END PORT
	END pin_565
	PIN pin_566
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 68.57868525896436 99.75 68.82868525896436 100 ;
		END PORT
	END pin_566
	PIN pin_567
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.25896414342651 99.75 68.50896414342651 100 ;
		END PORT
	END pin_567
	PIN pin_568
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 67.93924302788866 99.75 68.18924302788866 100 ;
		END PORT
	END pin_568
	PIN pin_569
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 67.61952191235082 99.75 67.86952191235082 100 ;
		END PORT
	END pin_569
	PIN pin_570
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.29980079681297 99.75 67.54980079681297 100 ;
		END PORT
	END pin_570
	PIN pin_571
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 66.98007968127513 99.75 67.23007968127513 100 ;
		END PORT
	END pin_571
	PIN pin_572
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 66.66035856573728 99.75 66.91035856573728 100 ;
		END PORT
	END pin_572
	PIN pin_573
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.34063745019944 99.75 66.59063745019944 100 ;
		END PORT
	END pin_573
	PIN pin_574
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.02091633466159 99.75 66.27091633466159 100 ;
		END PORT
	END pin_574
	PIN pin_575
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 65.70119521912375 99.75 65.95119521912375 100 ;
		END PORT
	END pin_575
	PIN pin_576
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 65.3814741035859 99.75 65.6314741035859 100 ;
		END PORT
	END pin_576
	PIN pin_577
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 65.06175298804806 99.75 65.31175298804806 100 ;
		END PORT
	END pin_577
	PIN pin_578
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.74203187251021 99.75 64.99203187251021 100 ;
		END PORT
	END pin_578
	PIN pin_579
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.42231075697237 99.75 64.67231075697237 100 ;
		END PORT
	END pin_579
	PIN pin_580
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.10258964143452 99.75 64.35258964143452 100 ;
		END PORT
	END pin_580
	PIN pin_581
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 63.782868525896674 99.75 64.03286852589667 100 ;
		END PORT
	END pin_581
	PIN pin_582
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.46314741035883 99.75 63.71314741035883 100 ;
		END PORT
	END pin_582
	PIN pin_583
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.14342629482098 99.75 63.39342629482098 100 ;
		END PORT
	END pin_583
	PIN pin_584
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 62.82370517928314 99.75 63.07370517928314 100 ;
		END PORT
	END pin_584
	PIN pin_585
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 62.50398406374529 99.75 62.75398406374529 100 ;
		END PORT
	END pin_585
	PIN pin_586
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 62.18426294820745 99.75 62.43426294820745 100 ;
		END PORT
	END pin_586
	PIN pin_587
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 61.8645418326696 99.75 62.1145418326696 100 ;
		END PORT
	END pin_587
	PIN pin_588
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 61.544820717131756 99.75 61.794820717131756 100 ;
		END PORT
	END pin_588
	PIN pin_589
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 61.22509960159391 99.75 61.47509960159391 100 ;
		END PORT
	END pin_589
	PIN pin_590
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 60.905378486056065 99.75 61.155378486056065 100 ;
		END PORT
	END pin_590
	PIN pin_591
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.58565737051822 99.75 60.83565737051822 100 ;
		END PORT
	END pin_591
	PIN pin_592
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.265936254980375 99.75 60.515936254980375 100 ;
		END PORT
	END pin_592
	PIN pin_593
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 59.94621513944253 99.75 60.19621513944253 100 ;
		END PORT
	END pin_593
	PIN pin_594
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 59.626494023904684 99.75 59.876494023904684 100 ;
		END PORT
	END pin_594
	PIN pin_595
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 59.30677290836684 99.75 59.55677290836684 100 ;
		END PORT
	END pin_595
	PIN pin_596
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.98705179282899 99.75 59.23705179282899 100 ;
		END PORT
	END pin_596
	PIN pin_597
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.66733067729115 99.75 58.91733067729115 100 ;
		END PORT
	END pin_597
	PIN pin_598
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.3476095617533 99.75 58.5976095617533 100 ;
		END PORT
	END pin_598
	PIN pin_599
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.02788844621546 99.75 58.27788844621546 100 ;
		END PORT
	END pin_599
	PIN pin_600
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 57.70816733067761 99.75 57.95816733067761 100 ;
		END PORT
	END pin_600
	PIN pin_601
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 57.388446215139766 99.75 57.638446215139766 100 ;
		END PORT
	END pin_601
	PIN pin_602
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 57.06872509960192 99.75 57.31872509960192 100 ;
		END PORT
	END pin_602
	PIN pin_603
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.749003984064075 99.75 56.999003984064075 100 ;
		END PORT
	END pin_603
	PIN pin_604
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.42928286852623 99.75 56.67928286852623 100 ;
		END PORT
	END pin_604
	PIN pin_605
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.109561752988384 99.75 56.359561752988384 100 ;
		END PORT
	END pin_605
	PIN pin_606
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 55.78984063745054 99.75 56.03984063745054 100 ;
		END PORT
	END pin_606
	PIN pin_607
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 55.47011952191269 99.75 55.72011952191269 100 ;
		END PORT
	END pin_607
	PIN pin_608
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.15039840637485 99.75 55.40039840637485 100 ;
		END PORT
	END pin_608
	PIN pin_609
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.830677290837 99.75 55.080677290837 100 ;
		END PORT
	END pin_609
	PIN pin_610
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.51095617529916 99.75 54.76095617529916 100 ;
		END PORT
	END pin_610
	PIN pin_611
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.19123505976131 99.75 54.44123505976131 100 ;
		END PORT
	END pin_611
	PIN pin_612
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 53.871513944223466 99.75 54.121513944223466 100 ;
		END PORT
	END pin_612
	PIN pin_613
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.55179282868562 99.75 53.80179282868562 100 ;
		END PORT
	END pin_613
	PIN pin_614
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 53.232071713147775 99.75 53.482071713147775 100 ;
		END PORT
	END pin_614
	PIN pin_615
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 52.91235059760993 99.75 53.16235059760993 100 ;
		END PORT
	END pin_615
	PIN pin_616
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 52.592629482072084 99.75 52.842629482072084 100 ;
		END PORT
	END pin_616
	PIN pin_617
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 52.27290836653424 99.75 52.52290836653424 100 ;
		END PORT
	END pin_617
	PIN pin_618
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.95318725099639 99.75 52.20318725099639 100 ;
		END PORT
	END pin_618
	PIN pin_619
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.63346613545855 99.75 51.88346613545855 100 ;
		END PORT
	END pin_619
	PIN pin_620
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 51.3137450199207 99.75 51.5637450199207 100 ;
		END PORT
	END pin_620
	PIN pin_621
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.99402390438286 99.75 51.24402390438286 100 ;
		END PORT
	END pin_621
	PIN pin_622
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 50.67430278884501 99.75 50.92430278884501 100 ;
		END PORT
	END pin_622
	PIN pin_623
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.354581673307166 99.75 50.604581673307166 100 ;
		END PORT
	END pin_623
	PIN pin_624
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.03486055776932 99.75 50.28486055776932 100 ;
		END PORT
	END pin_624
	PIN pin_625
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.715139442231475 99.75 49.965139442231475 100 ;
		END PORT
	END pin_625
	PIN pin_626
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.39541832669363 99.75 49.64541832669363 100 ;
		END PORT
	END pin_626
	PIN pin_627
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 49.075697211155784 99.75 49.325697211155784 100 ;
		END PORT
	END pin_627
	PIN pin_628
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 48.75597609561794 99.75 49.00597609561794 100 ;
		END PORT
	END pin_628
	PIN pin_629
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.43625498008009 99.75 48.68625498008009 100 ;
		END PORT
	END pin_629
	PIN pin_630
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 48.11653386454225 99.75 48.36653386454225 100 ;
		END PORT
	END pin_630
	PIN pin_631
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 47.7968127490044 99.75 48.0468127490044 100 ;
		END PORT
	END pin_631
	PIN pin_632
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.47709163346656 99.75 47.72709163346656 100 ;
		END PORT
	END pin_632
	PIN pin_633
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.15737051792871 99.75 47.40737051792871 100 ;
		END PORT
	END pin_633
	PIN pin_634
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.837649402390866 99.75 47.087649402390866 100 ;
		END PORT
	END pin_634
	PIN pin_635
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 46.51792828685302 99.75 46.76792828685302 100 ;
		END PORT
	END pin_635
	PIN pin_636
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.198207171315175 99.75 46.448207171315175 100 ;
		END PORT
	END pin_636
	PIN pin_637
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.87848605577733 99.75 46.12848605577733 100 ;
		END PORT
	END pin_637
	PIN pin_638
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.558764940239485 99.75 45.808764940239485 100 ;
		END PORT
	END pin_638
	PIN pin_639
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 45.23904382470164 99.75 45.48904382470164 100 ;
		END PORT
	END pin_639
	PIN pin_640
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 44.919322709163794 99.75 45.169322709163794 100 ;
		END PORT
	END pin_640
	PIN pin_641
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.59960159362595 99.75 44.84960159362595 100 ;
		END PORT
	END pin_641
	PIN pin_642
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 44.2798804780881 99.75 44.5298804780881 100 ;
		END PORT
	END pin_642
	PIN pin_643
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.96015936255026 99.75 44.21015936255026 100 ;
		END PORT
	END pin_643
	PIN pin_644
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 43.64043824701241 99.75 43.89043824701241 100 ;
		END PORT
	END pin_644
	PIN pin_645
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 43.32071713147457 99.75 43.57071713147457 100 ;
		END PORT
	END pin_645
	PIN pin_646
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 43.00099601593672 99.75 43.25099601593672 100 ;
		END PORT
	END pin_646
	PIN pin_647
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 42.681274900398876 99.75 42.931274900398876 100 ;
		END PORT
	END pin_647
	PIN pin_648
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.36155378486103 99.75 42.61155378486103 100 ;
		END PORT
	END pin_648
	PIN pin_649
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.041832669323185 99.75 42.291832669323185 100 ;
		END PORT
	END pin_649
	PIN pin_650
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 41.72211155378534 99.75 41.97211155378534 100 ;
		END PORT
	END pin_650
	PIN pin_651
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.402390438247494 99.75 41.652390438247494 100 ;
		END PORT
	END pin_651
	PIN pin_652
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.08266932270965 99.75 41.33266932270965 100 ;
		END PORT
	END pin_652
	PIN pin_653
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.7629482071718 99.75 41.0129482071718 100 ;
		END PORT
	END pin_653
	PIN pin_654
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 40.44322709163396 99.75 40.69322709163396 100 ;
		END PORT
	END pin_654
	PIN pin_655
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 40.12350597609611 99.75 40.37350597609611 100 ;
		END PORT
	END pin_655
	PIN pin_656
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 39.80378486055827 99.75 40.05378486055827 100 ;
		END PORT
	END pin_656
	PIN pin_657
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 39.48406374502042 99.75 39.73406374502042 100 ;
		END PORT
	END pin_657
	PIN pin_658
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 39.164342629482576 99.75 39.414342629482576 100 ;
		END PORT
	END pin_658
	PIN pin_659
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.84462151394473 99.75 39.09462151394473 100 ;
		END PORT
	END pin_659
	PIN pin_660
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 38.524900398406885 99.75 38.774900398406885 100 ;
		END PORT
	END pin_660
	PIN pin_661
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 38.20517928286904 99.75 38.45517928286904 100 ;
		END PORT
	END pin_661
	PIN pin_662
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.885458167331194 99.75 38.135458167331194 100 ;
		END PORT
	END pin_662
	PIN pin_663
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 37.56573705179335 99.75 37.81573705179335 100 ;
		END PORT
	END pin_663
	PIN pin_664
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 37.2460159362555 99.75 37.4960159362555 100 ;
		END PORT
	END pin_664
	PIN pin_665
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.92629482071766 99.75 37.17629482071766 100 ;
		END PORT
	END pin_665
	PIN pin_666
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 36.60657370517981 99.75 36.85657370517981 100 ;
		END PORT
	END pin_666
	PIN pin_667
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.28685258964197 99.75 36.53685258964197 100 ;
		END PORT
	END pin_667
	PIN pin_668
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 35.96713147410412 99.75 36.21713147410412 100 ;
		END PORT
	END pin_668
	PIN pin_669
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.647410358566276 99.75 35.897410358566276 100 ;
		END PORT
	END pin_669
	PIN pin_670
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 35.32768924302843 99.75 35.57768924302843 100 ;
		END PORT
	END pin_670
	PIN pin_671
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 35.007968127490585 99.75 35.257968127490585 100 ;
		END PORT
	END pin_671
	PIN pin_672
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.68824701195274 99.75 34.93824701195274 100 ;
		END PORT
	END pin_672
	PIN pin_673
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 34.368525896414894 99.75 34.618525896414894 100 ;
		END PORT
	END pin_673
	PIN pin_674
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.04880478087705 99.75 34.29880478087705 100 ;
		END PORT
	END pin_674
	PIN pin_675
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 33.7290836653392 99.75 33.9790836653392 100 ;
		END PORT
	END pin_675
	PIN pin_676
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.40936254980136 99.75 33.65936254980136 100 ;
		END PORT
	END pin_676
	PIN pin_677
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.08964143426351 99.75 33.33964143426351 100 ;
		END PORT
	END pin_677
	PIN pin_678
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.76992031872567 99.75 33.01992031872567 100 ;
		END PORT
	END pin_678
	PIN pin_679
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.45019920318782 99.75 32.70019920318782 100 ;
		END PORT
	END pin_679
	PIN pin_680
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.130478087649976 99.75 32.380478087649976 100 ;
		END PORT
	END pin_680
	PIN pin_681
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.81075697211213 99.75 32.06075697211213 100 ;
		END PORT
	END pin_681
	PIN pin_682
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.491035856574282 99.75 31.741035856574282 100 ;
		END PORT
	END pin_682
	PIN pin_683
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.171314741036433 99.75 31.421314741036433 100 ;
		END PORT
	END pin_683
	PIN pin_684
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 30.851593625498584 99.75 31.101593625498584 100 ;
		END PORT
	END pin_684
	PIN pin_685
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.531872509960735 99.75 30.781872509960735 100 ;
		END PORT
	END pin_685
	PIN pin_686
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.212151394422886 99.75 30.462151394422886 100 ;
		END PORT
	END pin_686
	PIN pin_687
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 29.892430278885037 99.75 30.142430278885037 100 ;
		END PORT
	END pin_687
	PIN pin_688
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 29.572709163347188 99.75 29.822709163347188 100 ;
		END PORT
	END pin_688
	PIN pin_689
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.25298804780934 99.75 29.50298804780934 100 ;
		END PORT
	END pin_689
	PIN pin_690
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 28.93326693227149 99.75 29.18326693227149 100 ;
		END PORT
	END pin_690
	PIN pin_691
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 28.61354581673364 99.75 28.86354581673364 100 ;
		END PORT
	END pin_691
	PIN pin_692
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.293824701195792 99.75 28.543824701195792 100 ;
		END PORT
	END pin_692
	PIN pin_693
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 27.974103585657943 99.75 28.224103585657943 100 ;
		END PORT
	END pin_693
	PIN pin_694
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.654382470120094 99.75 27.904382470120094 100 ;
		END PORT
	END pin_694
	PIN pin_695
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.334661354582245 99.75 27.584661354582245 100 ;
		END PORT
	END pin_695
	PIN pin_696
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 27.014940239044396 99.75 27.264940239044396 100 ;
		END PORT
	END pin_696
	PIN pin_697
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.695219123506547 99.75 26.945219123506547 100 ;
		END PORT
	END pin_697
	PIN pin_698
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.375498007968698 99.75 26.625498007968698 100 ;
		END PORT
	END pin_698
	PIN pin_699
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 26.05577689243085 99.75 26.30577689243085 100 ;
		END PORT
	END pin_699
	PIN pin_700
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 25.736055776893 99.75 25.986055776893 100 ;
		END PORT
	END pin_700
	PIN pin_701
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 25.41633466135515 99.75 25.66633466135515 100 ;
		END PORT
	END pin_701
	PIN pin_702
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 25.096613545817302 99.75 25.346613545817302 100 ;
		END PORT
	END pin_702
	PIN pin_703
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 24.776892430279453 99.75 25.026892430279453 100 ;
		END PORT
	END pin_703
	PIN pin_704
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.457171314741604 99.75 24.707171314741604 100 ;
		END PORT
	END pin_704
	PIN pin_705
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.137450199203755 99.75 24.387450199203755 100 ;
		END PORT
	END pin_705
	PIN pin_706
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 23.817729083665906 99.75 24.067729083665906 100 ;
		END PORT
	END pin_706
	PIN pin_707
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.498007968128057 99.75 23.748007968128057 100 ;
		END PORT
	END pin_707
	PIN pin_708
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.178286852590208 99.75 23.428286852590208 100 ;
		END PORT
	END pin_708
	PIN pin_709
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 22.85856573705236 99.75 23.10856573705236 100 ;
		END PORT
	END pin_709
	PIN pin_710
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 22.53884462151451 99.75 22.78884462151451 100 ;
		END PORT
	END pin_710
	PIN pin_711
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 22.21912350597666 99.75 22.46912350597666 100 ;
		END PORT
	END pin_711
	PIN pin_712
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 21.899402390438812 99.75 22.149402390438812 100 ;
		END PORT
	END pin_712
	PIN pin_713
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.579681274900963 99.75 21.829681274900963 100 ;
		END PORT
	END pin_713
	PIN pin_714
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 21.259960159363114 99.75 21.509960159363114 100 ;
		END PORT
	END pin_714
	PIN pin_715
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 20.940239043825265 99.75 21.190239043825265 100 ;
		END PORT
	END pin_715
	PIN pin_716
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.620517928287416 99.75 20.870517928287416 100 ;
		END PORT
	END pin_716
	PIN pin_717
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 20.300796812749567 99.75 20.550796812749567 100 ;
		END PORT
	END pin_717
	PIN pin_718
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 19.98107569721172 99.75 20.23107569721172 100 ;
		END PORT
	END pin_718
	PIN pin_719
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 19.66135458167387 99.75 19.91135458167387 100 ;
		END PORT
	END pin_719
	PIN pin_720
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 19.34163346613602 99.75 19.59163346613602 100 ;
		END PORT
	END pin_720
	PIN pin_721
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 19.02191235059817 99.75 19.27191235059817 100 ;
		END PORT
	END pin_721
	PIN pin_722
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 18.702191235060322 99.75 18.952191235060322 100 ;
		END PORT
	END pin_722
	PIN pin_723
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.382470119522473 99.75 18.632470119522473 100 ;
		END PORT
	END pin_723
	PIN pin_724
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 18.062749003984624 99.75 18.312749003984624 100 ;
		END PORT
	END pin_724
	PIN pin_725
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.743027888446775 99.75 17.993027888446775 100 ;
		END PORT
	END pin_725
	PIN pin_726
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 17.423306772908926 99.75 17.673306772908926 100 ;
		END PORT
	END pin_726
	PIN pin_727
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.103585657371077 99.75 17.353585657371077 100 ;
		END PORT
	END pin_727
	PIN pin_728
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.78386454183323 99.75 17.03386454183323 100 ;
		END PORT
	END pin_728
	PIN pin_729
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.46414342629538 99.75 16.71414342629538 100 ;
		END PORT
	END pin_729
	PIN pin_730
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.14442231075753 99.75 16.39442231075753 100 ;
		END PORT
	END pin_730
	PIN pin_731
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.824701195219681 99.75 16.07470119521968 100 ;
		END PORT
	END pin_731
	PIN pin_732
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 15.504980079681832 99.75 15.754980079681832 100 ;
		END PORT
	END pin_732
	PIN pin_733
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.185258964143983 99.75 15.435258964143983 100 ;
		END PORT
	END pin_733
	PIN pin_734
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.865537848606134 99.75 15.115537848606134 100 ;
		END PORT
	END pin_734
	PIN pin_735
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 14.545816733068285 99.75 14.795816733068285 100 ;
		END PORT
	END pin_735
	PIN pin_736
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 14.226095617530436 99.75 14.476095617530436 100 ;
		END PORT
	END pin_736
	PIN pin_737
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 13.906374501992588 99.75 14.156374501992588 100 ;
		END PORT
	END pin_737
	PIN pin_738
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 13.586653386454739 99.75 13.836653386454739 100 ;
		END PORT
	END pin_738
	PIN pin_739
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 13.26693227091689 99.75 13.51693227091689 100 ;
		END PORT
	END pin_739
	PIN pin_740
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 12.94721115537904 99.75 13.19721115537904 100 ;
		END PORT
	END pin_740
	PIN pin_741
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 12.627490039841192 99.75 12.877490039841192 100 ;
		END PORT
	END pin_741
	PIN pin_742
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 12.307768924303343 99.75 12.557768924303343 100 ;
		END PORT
	END pin_742
	PIN pin_743
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.988047808765494 99.75 12.238047808765494 100 ;
		END PORT
	END pin_743
	PIN pin_744
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 11.668326693227645 99.75 11.918326693227645 100 ;
		END PORT
	END pin_744
	PIN pin_745
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.348605577689796 99.75 11.598605577689796 100 ;
		END PORT
	END pin_745
	PIN pin_746
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.028884462151947 99.75 11.278884462151947 100 ;
		END PORT
	END pin_746
	PIN pin_747
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 10.709163346614098 99.75 10.959163346614098 100 ;
		END PORT
	END pin_747
	PIN pin_748
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 10.389442231076249 99.75 10.639442231076249 100 ;
		END PORT
	END pin_748
	PIN pin_749
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 10.0697211155384 99.75 10.3197211155384 100 ;
		END PORT
	END pin_749
	PIN pin_750
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 10.069721115537849 0 10.319721115537849 0.25 ;
		END PORT
	END pin_750
	PIN pin_751
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 10.389442231075698 0 10.639442231075698 0.25 ;
		END PORT
	END pin_751
	PIN pin_752
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 10.709163346613547 0 10.959163346613547 0.25 ;
		END PORT
	END pin_752
	PIN pin_753
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 11.028884462151396 0 11.278884462151396 0.25 ;
		END PORT
	END pin_753
	PIN pin_754
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.348605577689245 0 11.598605577689245 0.25 ;
		END PORT
	END pin_754
	PIN pin_755
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.668326693227094 0 11.918326693227094 0.25 ;
		END PORT
	END pin_755
	PIN pin_756
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.988047808764943 0 12.238047808764943 0.25 ;
		END PORT
	END pin_756
	PIN pin_757
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 12.307768924302792 0 12.557768924302792 0.25 ;
		END PORT
	END pin_757
	PIN pin_758
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 12.627490039840641 0 12.877490039840641 0.25 ;
		END PORT
	END pin_758
	PIN pin_759
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 12.94721115537849 0 13.19721115537849 0.25 ;
		END PORT
	END pin_759
	PIN pin_760
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 13.266932270916339 0 13.516932270916339 0.25 ;
		END PORT
	END pin_760
	PIN pin_761
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 13.586653386454188 0 13.836653386454188 0.25 ;
		END PORT
	END pin_761
	PIN pin_762
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 13.906374501992037 0 14.156374501992037 0.25 ;
		END PORT
	END pin_762
	PIN pin_763
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 14.226095617529886 0 14.476095617529886 0.25 ;
		END PORT
	END pin_763
	PIN pin_764
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 14.545816733067735 0 14.795816733067735 0.25 ;
		END PORT
	END pin_764
	PIN pin_765
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.865537848605584 0 15.115537848605584 0.25 ;
		END PORT
	END pin_765
	PIN pin_766
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.185258964143433 0 15.435258964143433 0.25 ;
		END PORT
	END pin_766
	PIN pin_767
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.504980079681282 0 15.754980079681282 0.25 ;
		END PORT
	END pin_767
	PIN pin_768
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.82470119521913 0 16.07470119521913 0.25 ;
		END PORT
	END pin_768
	PIN pin_769
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.14442231075698 0 16.39442231075698 0.25 ;
		END PORT
	END pin_769
	PIN pin_770
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.46414342629483 0 16.71414342629483 0.25 ;
		END PORT
	END pin_770
	PIN pin_771
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.783864541832678 0 17.033864541832678 0.25 ;
		END PORT
	END pin_771
	PIN pin_772
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 17.103585657370527 0 17.353585657370527 0.25 ;
		END PORT
	END pin_772
	PIN pin_773
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.423306772908376 0 17.673306772908376 0.25 ;
		END PORT
	END pin_773
	PIN pin_774
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 17.743027888446225 0 17.993027888446225 0.25 ;
		END PORT
	END pin_774
	PIN pin_775
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 18.062749003984074 0 18.312749003984074 0.25 ;
		END PORT
	END pin_775
	PIN pin_776
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.382470119521923 0 18.632470119521923 0.25 ;
		END PORT
	END pin_776
	PIN pin_777
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 18.70219123505977 0 18.95219123505977 0.25 ;
		END PORT
	END pin_777
	PIN pin_778
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.02191235059762 0 19.27191235059762 0.25 ;
		END PORT
	END pin_778
	PIN pin_779
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.34163346613547 0 19.59163346613547 0.25 ;
		END PORT
	END pin_779
	PIN pin_780
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.66135458167332 0 19.91135458167332 0.25 ;
		END PORT
	END pin_780
	PIN pin_781
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.981075697211168 0 20.231075697211168 0.25 ;
		END PORT
	END pin_781
	PIN pin_782
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.300796812749017 0 20.550796812749017 0.25 ;
		END PORT
	END pin_782
	PIN pin_783
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 20.620517928286866 0 20.870517928286866 0.25 ;
		END PORT
	END pin_783
	PIN pin_784
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.940239043824715 0 21.190239043824715 0.25 ;
		END PORT
	END pin_784
	PIN pin_785
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.259960159362564 0 21.509960159362564 0.25 ;
		END PORT
	END pin_785
	PIN pin_786
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 21.579681274900413 0 21.829681274900413 0.25 ;
		END PORT
	END pin_786
	PIN pin_787
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.89940239043826 0 22.14940239043826 0.25 ;
		END PORT
	END pin_787
	PIN pin_788
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 22.21912350597611 0 22.46912350597611 0.25 ;
		END PORT
	END pin_788
	PIN pin_789
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 22.53884462151396 0 22.78884462151396 0.25 ;
		END PORT
	END pin_789
	PIN pin_790
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.85856573705181 0 23.10856573705181 0.25 ;
		END PORT
	END pin_790
	PIN pin_791
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 23.178286852589657 0 23.428286852589657 0.25 ;
		END PORT
	END pin_791
	PIN pin_792
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 23.498007968127506 0 23.748007968127506 0.25 ;
		END PORT
	END pin_792
	PIN pin_793
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.817729083665355 0 24.067729083665355 0.25 ;
		END PORT
	END pin_793
	PIN pin_794
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.137450199203204 0 24.387450199203204 0.25 ;
		END PORT
	END pin_794
	PIN pin_795
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.457171314741053 0 24.707171314741053 0.25 ;
		END PORT
	END pin_795
	PIN pin_796
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 24.776892430278902 0 25.026892430278902 0.25 ;
		END PORT
	END pin_796
	PIN pin_797
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 25.09661354581675 0 25.34661354581675 0.25 ;
		END PORT
	END pin_797
	PIN pin_798
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 25.4163346613546 0 25.6663346613546 0.25 ;
		END PORT
	END pin_798
	PIN pin_799
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 25.73605577689245 0 25.98605577689245 0.25 ;
		END PORT
	END pin_799
	PIN pin_800
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.0557768924303 0 26.3057768924303 0.25 ;
		END PORT
	END pin_800
	PIN pin_801
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 26.375498007968147 0 26.625498007968147 0.25 ;
		END PORT
	END pin_801
	PIN pin_802
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 26.695219123505996 0 26.945219123505996 0.25 ;
		END PORT
	END pin_802
	PIN pin_803
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.014940239043845 0 27.264940239043845 0.25 ;
		END PORT
	END pin_803
	PIN pin_804
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 27.334661354581694 0 27.584661354581694 0.25 ;
		END PORT
	END pin_804
	PIN pin_805
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.654382470119543 0 27.904382470119543 0.25 ;
		END PORT
	END pin_805
	PIN pin_806
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.974103585657392 0 28.224103585657392 0.25 ;
		END PORT
	END pin_806
	PIN pin_807
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 28.29382470119524 0 28.54382470119524 0.25 ;
		END PORT
	END pin_807
	PIN pin_808
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 28.61354581673309 0 28.86354581673309 0.25 ;
		END PORT
	END pin_808
	PIN pin_809
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.93326693227094 0 29.18326693227094 0.25 ;
		END PORT
	END pin_809
	PIN pin_810
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.25298804780879 0 29.50298804780879 0.25 ;
		END PORT
	END pin_810
	PIN pin_811
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 29.572709163346637 0 29.822709163346637 0.25 ;
		END PORT
	END pin_811
	PIN pin_812
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.892430278884486 0 30.142430278884486 0.25 ;
		END PORT
	END pin_812
	PIN pin_813
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.212151394422335 0 30.462151394422335 0.25 ;
		END PORT
	END pin_813
	PIN pin_814
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 30.531872509960184 0 30.781872509960184 0.25 ;
		END PORT
	END pin_814
	PIN pin_815
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.851593625498033 0 31.101593625498033 0.25 ;
		END PORT
	END pin_815
	PIN pin_816
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 31.171314741035882 0 31.421314741035882 0.25 ;
		END PORT
	END pin_816
	PIN pin_817
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.49103585657373 0 31.74103585657373 0.25 ;
		END PORT
	END pin_817
	PIN pin_818
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.81075697211158 0 32.06075697211158 0.25 ;
		END PORT
	END pin_818
	PIN pin_819
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 32.13047808764942 0 32.38047808764942 0.25 ;
		END PORT
	END pin_819
	PIN pin_820
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.45019920318727 0 32.70019920318727 0.25 ;
		END PORT
	END pin_820
	PIN pin_821
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 32.76992031872511 0 33.01992031872511 0.25 ;
		END PORT
	END pin_821
	PIN pin_822
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 33.08964143426296 0 33.33964143426296 0.25 ;
		END PORT
	END pin_822
	PIN pin_823
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 33.409362549800804 0 33.659362549800804 0.25 ;
		END PORT
	END pin_823
	PIN pin_824
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.72908366533865 0 33.97908366533865 0.25 ;
		END PORT
	END pin_824
	PIN pin_825
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 34.048804780876495 0 34.298804780876495 0.25 ;
		END PORT
	END pin_825
	PIN pin_826
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 34.36852589641434 0 34.61852589641434 0.25 ;
		END PORT
	END pin_826
	PIN pin_827
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 34.688247011952186 0 34.938247011952186 0.25 ;
		END PORT
	END pin_827
	PIN pin_828
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 35.00796812749003 0 35.25796812749003 0.25 ;
		END PORT
	END pin_828
	PIN pin_829
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.327689243027876 0 35.577689243027876 0.25 ;
		END PORT
	END pin_829
	PIN pin_830
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.64741035856572 0 35.89741035856572 0.25 ;
		END PORT
	END pin_830
	PIN pin_831
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 35.96713147410357 0 36.21713147410357 0.25 ;
		END PORT
	END pin_831
	PIN pin_832
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 36.28685258964141 0 36.53685258964141 0.25 ;
		END PORT
	END pin_832
	PIN pin_833
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 36.60657370517926 0 36.85657370517926 0.25 ;
		END PORT
	END pin_833
	PIN pin_834
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 36.926294820717104 0 37.176294820717104 0.25 ;
		END PORT
	END pin_834
	PIN pin_835
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 37.24601593625495 0 37.49601593625495 0.25 ;
		END PORT
	END pin_835
	PIN pin_836
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.565737051792794 0 37.815737051792794 0.25 ;
		END PORT
	END pin_836
	PIN pin_837
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 37.88545816733064 0 38.13545816733064 0.25 ;
		END PORT
	END pin_837
	PIN pin_838
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 38.205179282868485 0 38.455179282868485 0.25 ;
		END PORT
	END pin_838
	PIN pin_839
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 38.52490039840633 0 38.77490039840633 0.25 ;
		END PORT
	END pin_839
	PIN pin_840
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.844621513944176 0 39.094621513944176 0.25 ;
		END PORT
	END pin_840
	PIN pin_841
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 39.16434262948202 0 39.41434262948202 0.25 ;
		END PORT
	END pin_841
	PIN pin_842
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 39.48406374501987 0 39.73406374501987 0.25 ;
		END PORT
	END pin_842
	PIN pin_843
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 39.80378486055771 0 40.05378486055771 0.25 ;
		END PORT
	END pin_843
	PIN pin_844
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.12350597609556 0 40.37350597609556 0.25 ;
		END PORT
	END pin_844
	PIN pin_845
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.4432270916334 0 40.6932270916334 0.25 ;
		END PORT
	END pin_845
	PIN pin_846
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.76294820717125 0 41.01294820717125 0.25 ;
		END PORT
	END pin_846
	PIN pin_847
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.082669322709094 0 41.332669322709094 0.25 ;
		END PORT
	END pin_847
	PIN pin_848
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 41.40239043824694 0 41.65239043824694 0.25 ;
		END PORT
	END pin_848
	PIN pin_849
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 41.722111553784785 0 41.972111553784785 0.25 ;
		END PORT
	END pin_849
	PIN pin_850
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 42.04183266932263 0 42.29183266932263 0.25 ;
		END PORT
	END pin_850
	PIN pin_851
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 42.361553784860476 0 42.611553784860476 0.25 ;
		END PORT
	END pin_851
	PIN pin_852
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.68127490039832 0 42.93127490039832 0.25 ;
		END PORT
	END pin_852
	PIN pin_853
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 43.00099601593617 0 43.25099601593617 0.25 ;
		END PORT
	END pin_853
	PIN pin_854
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 43.32071713147401 0 43.57071713147401 0.25 ;
		END PORT
	END pin_854
	PIN pin_855
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.64043824701186 0 43.89043824701186 0.25 ;
		END PORT
	END pin_855
	PIN pin_856
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.9601593625497 0 44.2101593625497 0.25 ;
		END PORT
	END pin_856
	PIN pin_857
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.27988047808755 0 44.52988047808755 0.25 ;
		END PORT
	END pin_857
	PIN pin_858
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.599601593625394 0 44.849601593625394 0.25 ;
		END PORT
	END pin_858
	PIN pin_859
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 44.91932270916324 0 45.16932270916324 0.25 ;
		END PORT
	END pin_859
	PIN pin_860
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 45.239043824701085 0 45.489043824701085 0.25 ;
		END PORT
	END pin_860
	PIN pin_861
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.55876494023893 0 45.80876494023893 0.25 ;
		END PORT
	END pin_861
	PIN pin_862
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.878486055776776 0 46.128486055776776 0.25 ;
		END PORT
	END pin_862
	PIN pin_863
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 46.19820717131462 0 46.44820717131462 0.25 ;
		END PORT
	END pin_863
	PIN pin_864
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.51792828685247 0 46.76792828685247 0.25 ;
		END PORT
	END pin_864
	PIN pin_865
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.83764940239031 0 47.08764940239031 0.25 ;
		END PORT
	END pin_865
	PIN pin_866
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.15737051792816 0 47.40737051792816 0.25 ;
		END PORT
	END pin_866
	PIN pin_867
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.477091633466 0 47.727091633466 0.25 ;
		END PORT
	END pin_867
	PIN pin_868
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.79681274900385 0 48.04681274900385 0.25 ;
		END PORT
	END pin_868
	PIN pin_869
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.116533864541694 0 48.366533864541694 0.25 ;
		END PORT
	END pin_869
	PIN pin_870
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 48.43625498007954 0 48.68625498007954 0.25 ;
		END PORT
	END pin_870
	PIN pin_871
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.755976095617385 0 49.005976095617385 0.25 ;
		END PORT
	END pin_871
	PIN pin_872
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 49.07569721115523 0 49.32569721115523 0.25 ;
		END PORT
	END pin_872
	PIN pin_873
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.395418326693076 0 49.645418326693076 0.25 ;
		END PORT
	END pin_873
	PIN pin_874
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 49.71513944223092 0 49.96513944223092 0.25 ;
		END PORT
	END pin_874
	PIN pin_875
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.034860557768766 0 50.284860557768766 0.25 ;
		END PORT
	END pin_875
	PIN pin_876
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 50.35458167330661 0 50.60458167330661 0.25 ;
		END PORT
	END pin_876
	PIN pin_877
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.67430278884446 0 50.92430278884446 0.25 ;
		END PORT
	END pin_877
	PIN pin_878
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.9940239043823 0 51.2440239043823 0.25 ;
		END PORT
	END pin_878
	PIN pin_879
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.31374501992015 0 51.56374501992015 0.25 ;
		END PORT
	END pin_879
	PIN pin_880
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 51.633466135457994 0 51.883466135457994 0.25 ;
		END PORT
	END pin_880
	PIN pin_881
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 51.95318725099584 0 52.20318725099584 0.25 ;
		END PORT
	END pin_881
	PIN pin_882
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 52.272908366533684 0 52.522908366533684 0.25 ;
		END PORT
	END pin_882
	PIN pin_883
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 52.59262948207153 0 52.84262948207153 0.25 ;
		END PORT
	END pin_883
	PIN pin_884
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 52.912350597609375 0 53.162350597609375 0.25 ;
		END PORT
	END pin_884
	PIN pin_885
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 53.23207171314722 0 53.48207171314722 0.25 ;
		END PORT
	END pin_885
	PIN pin_886
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 53.551792828685066 0 53.801792828685066 0.25 ;
		END PORT
	END pin_886
	PIN pin_887
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.87151394422291 0 54.12151394422291 0.25 ;
		END PORT
	END pin_887
	PIN pin_888
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 54.19123505976076 0 54.44123505976076 0.25 ;
		END PORT
	END pin_888
	PIN pin_889
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 54.5109561752986 0 54.7609561752986 0.25 ;
		END PORT
	END pin_889
	PIN pin_890
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.83067729083645 0 55.08067729083645 0.25 ;
		END PORT
	END pin_890
	PIN pin_891
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.15039840637429 0 55.40039840637429 0.25 ;
		END PORT
	END pin_891
	PIN pin_892
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 55.47011952191214 0 55.72011952191214 0.25 ;
		END PORT
	END pin_892
	PIN pin_893
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.789840637449984 0 56.039840637449984 0.25 ;
		END PORT
	END pin_893
	PIN pin_894
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.10956175298783 0 56.35956175298783 0.25 ;
		END PORT
	END pin_894
	PIN pin_895
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.429282868525675 0 56.679282868525675 0.25 ;
		END PORT
	END pin_895
	PIN pin_896
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.74900398406352 0 56.99900398406352 0.25 ;
		END PORT
	END pin_896
	PIN pin_897
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.068725099601366 0 57.318725099601366 0.25 ;
		END PORT
	END pin_897
	PIN pin_898
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 57.38844621513921 0 57.63844621513921 0.25 ;
		END PORT
	END pin_898
	PIN pin_899
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.70816733067706 0 57.95816733067706 0.25 ;
		END PORT
	END pin_899
	PIN pin_900
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.0278884462149 0 58.2778884462149 0.25 ;
		END PORT
	END pin_900
	PIN pin_901
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.34760956175275 0 58.59760956175275 0.25 ;
		END PORT
	END pin_901
	PIN pin_902
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.66733067729059 0 58.91733067729059 0.25 ;
		END PORT
	END pin_902
	PIN pin_903
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.98705179282844 0 59.23705179282844 0.25 ;
		END PORT
	END pin_903
	PIN pin_904
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 59.306772908366284 0 59.556772908366284 0.25 ;
		END PORT
	END pin_904
	PIN pin_905
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 59.62649402390413 0 59.87649402390413 0.25 ;
		END PORT
	END pin_905
	PIN pin_906
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 59.946215139441975 0 60.196215139441975 0.25 ;
		END PORT
	END pin_906
	PIN pin_907
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 60.26593625497982 0 60.51593625497982 0.25 ;
		END PORT
	END pin_907
	PIN pin_908
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 60.585657370517666 0 60.835657370517666 0.25 ;
		END PORT
	END pin_908
	PIN pin_909
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.90537848605551 0 61.15537848605551 0.25 ;
		END PORT
	END pin_909
	PIN pin_910
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 61.22509960159336 0 61.47509960159336 0.25 ;
		END PORT
	END pin_910
	PIN pin_911
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 61.5448207171312 0 61.7948207171312 0.25 ;
		END PORT
	END pin_911
	PIN pin_912
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 61.86454183266905 0 62.11454183266905 0.25 ;
		END PORT
	END pin_912
	PIN pin_913
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.18426294820689 0 62.43426294820689 0.25 ;
		END PORT
	END pin_913
	PIN pin_914
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 62.50398406374474 0 62.75398406374474 0.25 ;
		END PORT
	END pin_914
	PIN pin_915
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 62.823705179282584 0 63.073705179282584 0.25 ;
		END PORT
	END pin_915
	PIN pin_916
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.14342629482043 0 63.39342629482043 0.25 ;
		END PORT
	END pin_916
	PIN pin_917
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.463147410358275 0 63.713147410358275 0.25 ;
		END PORT
	END pin_917
	PIN pin_918
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.78286852589612 0 64.03286852589612 0.25 ;
		END PORT
	END pin_918
	PIN pin_919
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.10258964143397 0 64.35258964143397 0.25 ;
		END PORT
	END pin_919
	PIN pin_920
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.42231075697181 0 64.67231075697181 0.25 ;
		END PORT
	END pin_920
	PIN pin_921
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 64.74203187250966 0 64.99203187250966 0.25 ;
		END PORT
	END pin_921
	PIN pin_922
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.0617529880475 0 65.3117529880475 0.25 ;
		END PORT
	END pin_922
	PIN pin_923
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.38147410358535 0 65.63147410358535 0.25 ;
		END PORT
	END pin_923
	PIN pin_924
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.70119521912319 0 65.95119521912319 0.25 ;
		END PORT
	END pin_924
	PIN pin_925
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 66.02091633466104 0 66.27091633466104 0.25 ;
		END PORT
	END pin_925
	PIN pin_926
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 66.34063745019888 0 66.59063745019888 0.25 ;
		END PORT
	END pin_926
	PIN pin_927
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.66035856573673 0 66.91035856573673 0.25 ;
		END PORT
	END pin_927
	PIN pin_928
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.98007968127457 0 67.23007968127457 0.25 ;
		END PORT
	END pin_928
	PIN pin_929
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 67.29980079681242 0 67.54980079681242 0.25 ;
		END PORT
	END pin_929
	PIN pin_930
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 67.61952191235027 0 67.86952191235027 0.25 ;
		END PORT
	END pin_930
	PIN pin_931
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.93924302788811 0 68.18924302788811 0.25 ;
		END PORT
	END pin_931
	PIN pin_932
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 68.25896414342596 0 68.50896414342596 0.25 ;
		END PORT
	END pin_932
	PIN pin_933
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.5786852589638 0 68.8286852589638 0.25 ;
		END PORT
	END pin_933
	PIN pin_934
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 68.89840637450165 0 69.14840637450165 0.25 ;
		END PORT
	END pin_934
	PIN pin_935
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 69.21812749003949 0 69.46812749003949 0.25 ;
		END PORT
	END pin_935
	PIN pin_936
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 69.53784860557734 0 69.78784860557734 0.25 ;
		END PORT
	END pin_936
	PIN pin_937
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 69.85756972111518 0 70.10756972111518 0.25 ;
		END PORT
	END pin_937
	PIN pin_938
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 70.17729083665303 0 70.42729083665303 0.25 ;
		END PORT
	END pin_938
	PIN pin_939
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.49701195219087 0 70.74701195219087 0.25 ;
		END PORT
	END pin_939
	PIN pin_940
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 70.81673306772872 0 71.06673306772872 0.25 ;
		END PORT
	END pin_940
	PIN pin_941
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 71.13645418326657 0 71.38645418326657 0.25 ;
		END PORT
	END pin_941
	PIN pin_942
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 71.45617529880441 0 71.70617529880441 0.25 ;
		END PORT
	END pin_942
	PIN pin_943
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 71.77589641434226 0 72.02589641434226 0.25 ;
		END PORT
	END pin_943
	PIN pin_944
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 72.0956175298801 0 72.3456175298801 0.25 ;
		END PORT
	END pin_944
	PIN pin_945
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 72.41533864541795 0 72.66533864541795 0.25 ;
		END PORT
	END pin_945
	PIN pin_946
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 72.73505976095579 0 72.98505976095579 0.25 ;
		END PORT
	END pin_946
	PIN pin_947
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 73.05478087649364 0 73.30478087649364 0.25 ;
		END PORT
	END pin_947
	PIN pin_948
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.37450199203148 0 73.62450199203148 0.25 ;
		END PORT
	END pin_948
	PIN pin_949
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.69422310756933 0 73.94422310756933 0.25 ;
		END PORT
	END pin_949
	PIN pin_950
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 74.01394422310717 0 74.26394422310717 0.25 ;
		END PORT
	END pin_950
	PIN pin_951
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.33366533864502 0 74.58366533864502 0.25 ;
		END PORT
	END pin_951
	PIN pin_952
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.65338645418286 0 74.90338645418286 0.25 ;
		END PORT
	END pin_952
	PIN pin_953
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 74.97310756972071 0 75.22310756972071 0.25 ;
		END PORT
	END pin_953
	PIN pin_954
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.29282868525856 0 75.54282868525856 0.25 ;
		END PORT
	END pin_954
	PIN pin_955
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 75.6125498007964 0 75.8625498007964 0.25 ;
		END PORT
	END pin_955
	PIN pin_956
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 75.93227091633425 0 76.18227091633425 0.25 ;
		END PORT
	END pin_956
	PIN pin_957
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 76.25199203187209 0 76.50199203187209 0.25 ;
		END PORT
	END pin_957
	PIN pin_958
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 76.57171314740994 0 76.82171314740994 0.25 ;
		END PORT
	END pin_958
	PIN pin_959
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 76.89143426294778 0 77.14143426294778 0.25 ;
		END PORT
	END pin_959
	PIN pin_960
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.21115537848563 0 77.46115537848563 0.25 ;
		END PORT
	END pin_960
	PIN pin_961
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 77.53087649402347 0 77.78087649402347 0.25 ;
		END PORT
	END pin_961
	PIN pin_962
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 77.85059760956132 0 78.10059760956132 0.25 ;
		END PORT
	END pin_962
	PIN pin_963
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 78.17031872509916 0 78.42031872509916 0.25 ;
		END PORT
	END pin_963
	PIN pin_964
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 78.49003984063701 0 78.74003984063701 0.25 ;
		END PORT
	END pin_964
	PIN pin_965
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 78.80976095617486 0 79.05976095617486 0.25 ;
		END PORT
	END pin_965
	PIN pin_966
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.1294820717127 0 79.3794820717127 0.25 ;
		END PORT
	END pin_966
	PIN pin_967
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.44920318725055 0 79.69920318725055 0.25 ;
		END PORT
	END pin_967
	PIN pin_968
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.76892430278839 0 80.01892430278839 0.25 ;
		END PORT
	END pin_968
	PIN pin_969
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 80.08864541832624 0 80.33864541832624 0.25 ;
		END PORT
	END pin_969
	PIN pin_970
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.40836653386408 0 80.65836653386408 0.25 ;
		END PORT
	END pin_970
	PIN pin_971
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 80.72808764940193 0 80.97808764940193 0.25 ;
		END PORT
	END pin_971
	PIN pin_972
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.04780876493977 0 81.29780876493977 0.25 ;
		END PORT
	END pin_972
	PIN pin_973
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.36752988047762 0 81.61752988047762 0.25 ;
		END PORT
	END pin_973
	PIN pin_974
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.68725099601546 0 81.93725099601546 0.25 ;
		END PORT
	END pin_974
	PIN pin_975
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.00697211155331 0 82.25697211155331 0.25 ;
		END PORT
	END pin_975
	PIN pin_976
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.32669322709116 0 82.57669322709116 0.25 ;
		END PORT
	END pin_976
	PIN pin_977
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.646414342629 0 82.896414342629 0.25 ;
		END PORT
	END pin_977
	PIN pin_978
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.96613545816685 0 83.21613545816685 0.25 ;
		END PORT
	END pin_978
	PIN pin_979
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.28585657370469 0 83.53585657370469 0.25 ;
		END PORT
	END pin_979
	PIN pin_980
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 83.60557768924254 0 83.85557768924254 0.25 ;
		END PORT
	END pin_980
	PIN pin_981
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.92529880478038 0 84.17529880478038 0.25 ;
		END PORT
	END pin_981
	PIN pin_982
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 84.24501992031823 0 84.49501992031823 0.25 ;
		END PORT
	END pin_982
	PIN pin_983
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 84.56474103585607 0 84.81474103585607 0.25 ;
		END PORT
	END pin_983
	PIN pin_984
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 84.88446215139392 0 85.13446215139392 0.25 ;
		END PORT
	END pin_984
	PIN pin_985
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 85.20418326693176 0 85.45418326693176 0.25 ;
		END PORT
	END pin_985
	PIN pin_986
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 85.52390438246961 0 85.77390438246961 0.25 ;
		END PORT
	END pin_986
	PIN pin_987
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.84362549800746 0 86.09362549800746 0.25 ;
		END PORT
	END pin_987
	PIN pin_988
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 86.1633466135453 0 86.4133466135453 0.25 ;
		END PORT
	END pin_988
	PIN pin_989
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.48306772908315 0 86.73306772908315 0.25 ;
		END PORT
	END pin_989
	PIN pin_990
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 86.80278884462099 0 87.05278884462099 0.25 ;
		END PORT
	END pin_990
	PIN pin_991
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 87.12250996015884 0 87.37250996015884 0.25 ;
		END PORT
	END pin_991
	PIN pin_992
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.44223107569668 0 87.69223107569668 0.25 ;
		END PORT
	END pin_992
	PIN pin_993
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.76195219123453 0 88.01195219123453 0.25 ;
		END PORT
	END pin_993
	PIN pin_994
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 88.08167330677237 0 88.33167330677237 0.25 ;
		END PORT
	END pin_994
	PIN pin_995
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 88.40139442231022 0 88.65139442231022 0.25 ;
		END PORT
	END pin_995
	PIN pin_996
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 88.72111553784806 0 88.97111553784806 0.25 ;
		END PORT
	END pin_996
	PIN pin_997
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.04083665338591 0 89.29083665338591 0.25 ;
		END PORT
	END pin_997
	PIN pin_998
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 89.36055776892375 0 89.61055776892375 0.25 ;
		END PORT
	END pin_998
	PIN pin_999
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.6802788844616 0 89.9302788844616 0.25 ;
		END PORT
	END pin_999
END MACRO
MACRO cell_1
	SIZE 100 BY 100 ;
	PIN pin_0
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 89.68027888446215 0.25 89.93027888446215 ;
		END PORT
	END pin_0
	PIN pin_1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 89.36055776892431 0.25 89.61055776892431 ;
		END PORT
	END pin_1
	PIN pin_2
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 89.04083665338646 0.25 89.29083665338646 ;
		END PORT
	END pin_2
	PIN pin_3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 88.72111553784862 0.25 88.97111553784862 ;
		END PORT
	END pin_3
	PIN pin_4
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 88.40139442231077 0.25 88.65139442231077 ;
		END PORT
	END pin_4
	PIN pin_5
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 88.08167330677293 0.25 88.33167330677293 ;
		END PORT
	END pin_5
	PIN pin_6
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 87.76195219123508 0.25 88.01195219123508 ;
		END PORT
	END pin_6
	PIN pin_7
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 87.44223107569724 0.25 87.69223107569724 ;
		END PORT
	END pin_7
	PIN pin_8
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 87.12250996015939 0.25 87.37250996015939 ;
		END PORT
	END pin_8
	PIN pin_9
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 86.80278884462155 0.25 87.05278884462155 ;
		END PORT
	END pin_9
	PIN pin_10
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 86.4830677290837 0.25 86.7330677290837 ;
		END PORT
	END pin_10
	PIN pin_11
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 86.16334661354585 0.25 86.41334661354585 ;
		END PORT
	END pin_11
	PIN pin_12
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 85.84362549800801 0.25 86.09362549800801 ;
		END PORT
	END pin_12
	PIN pin_13
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 85.52390438247016 0.25 85.77390438247016 ;
		END PORT
	END pin_13
	PIN pin_14
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 85.20418326693232 0.25 85.45418326693232 ;
		END PORT
	END pin_14
	PIN pin_15
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 84.88446215139447 0.25 85.13446215139447 ;
		END PORT
	END pin_15
	PIN pin_16
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 84.56474103585663 0.25 84.81474103585663 ;
		END PORT
	END pin_16
	PIN pin_17
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 84.24501992031878 0.25 84.49501992031878 ;
		END PORT
	END pin_17
	PIN pin_18
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 83.92529880478094 0.25 84.17529880478094 ;
		END PORT
	END pin_18
	PIN pin_19
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 83.60557768924309 0.25 83.85557768924309 ;
		END PORT
	END pin_19
	PIN pin_20
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 83.28585657370525 0.25 83.53585657370525 ;
		END PORT
	END pin_20
	PIN pin_21
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 82.9661354581674 0.25 83.2161354581674 ;
		END PORT
	END pin_21
	PIN pin_22
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 82.64641434262955 0.25 82.89641434262955 ;
		END PORT
	END pin_22
	PIN pin_23
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 82.32669322709171 0.25 82.57669322709171 ;
		END PORT
	END pin_23
	PIN pin_24
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 82.00697211155386 0.25 82.25697211155386 ;
		END PORT
	END pin_24
	PIN pin_25
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 81.68725099601602 0.25 81.93725099601602 ;
		END PORT
	END pin_25
	PIN pin_26
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 81.36752988047817 0.25 81.61752988047817 ;
		END PORT
	END pin_26
	PIN pin_27
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 81.04780876494033 0.25 81.29780876494033 ;
		END PORT
	END pin_27
	PIN pin_28
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 80.72808764940248 0.25 80.97808764940248 ;
		END PORT
	END pin_28
	PIN pin_29
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 80.40836653386464 0.25 80.65836653386464 ;
		END PORT
	END pin_29
	PIN pin_30
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 80.08864541832679 0.25 80.33864541832679 ;
		END PORT
	END pin_30
	PIN pin_31
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 79.76892430278895 0.25 80.01892430278895 ;
		END PORT
	END pin_31
	PIN pin_32
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 79.4492031872511 0.25 79.6992031872511 ;
		END PORT
	END pin_32
	PIN pin_33
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 79.12948207171326 0.25 79.37948207171326 ;
		END PORT
	END pin_33
	PIN pin_34
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 78.80976095617541 0.25 79.05976095617541 ;
		END PORT
	END pin_34
	PIN pin_35
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 78.49003984063756 0.25 78.74003984063756 ;
		END PORT
	END pin_35
	PIN pin_36
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 78.17031872509972 0.25 78.42031872509972 ;
		END PORT
	END pin_36
	PIN pin_37
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 77.85059760956187 0.25 78.10059760956187 ;
		END PORT
	END pin_37
	PIN pin_38
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 77.53087649402403 0.25 77.78087649402403 ;
		END PORT
	END pin_38
	PIN pin_39
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 77.21115537848618 0.25 77.46115537848618 ;
		END PORT
	END pin_39
	PIN pin_40
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 76.89143426294834 0.25 77.14143426294834 ;
		END PORT
	END pin_40
	PIN pin_41
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 76.57171314741049 0.25 76.82171314741049 ;
		END PORT
	END pin_41
	PIN pin_42
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 76.25199203187265 0.25 76.50199203187265 ;
		END PORT
	END pin_42
	PIN pin_43
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 75.9322709163348 0.25 76.1822709163348 ;
		END PORT
	END pin_43
	PIN pin_44
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 75.61254980079696 0.25 75.86254980079696 ;
		END PORT
	END pin_44
	PIN pin_45
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 75.29282868525911 0.25 75.54282868525911 ;
		END PORT
	END pin_45
	PIN pin_46
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 74.97310756972126 0.25 75.22310756972126 ;
		END PORT
	END pin_46
	PIN pin_47
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 74.65338645418342 0.25 74.90338645418342 ;
		END PORT
	END pin_47
	PIN pin_48
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 74.33366533864557 0.25 74.58366533864557 ;
		END PORT
	END pin_48
	PIN pin_49
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 74.01394422310773 0.25 74.26394422310773 ;
		END PORT
	END pin_49
	PIN pin_50
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 73.69422310756988 0.25 73.94422310756988 ;
		END PORT
	END pin_50
	PIN pin_51
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 73.37450199203204 0.25 73.62450199203204 ;
		END PORT
	END pin_51
	PIN pin_52
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 73.05478087649419 0.25 73.30478087649419 ;
		END PORT
	END pin_52
	PIN pin_53
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 72.73505976095635 0.25 72.98505976095635 ;
		END PORT
	END pin_53
	PIN pin_54
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 72.4153386454185 0.25 72.6653386454185 ;
		END PORT
	END pin_54
	PIN pin_55
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 72.09561752988066 0.25 72.34561752988066 ;
		END PORT
	END pin_55
	PIN pin_56
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 71.77589641434281 0.25 72.02589641434281 ;
		END PORT
	END pin_56
	PIN pin_57
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 71.45617529880496 0.25 71.70617529880496 ;
		END PORT
	END pin_57
	PIN pin_58
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 71.13645418326712 0.25 71.38645418326712 ;
		END PORT
	END pin_58
	PIN pin_59
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 70.81673306772927 0.25 71.06673306772927 ;
		END PORT
	END pin_59
	PIN pin_60
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 70.49701195219143 0.25 70.74701195219143 ;
		END PORT
	END pin_60
	PIN pin_61
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 70.17729083665358 0.25 70.42729083665358 ;
		END PORT
	END pin_61
	PIN pin_62
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 69.85756972111574 0.25 70.10756972111574 ;
		END PORT
	END pin_62
	PIN pin_63
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 69.53784860557789 0.25 69.78784860557789 ;
		END PORT
	END pin_63
	PIN pin_64
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 69.21812749004005 0.25 69.46812749004005 ;
		END PORT
	END pin_64
	PIN pin_65
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 68.8984063745022 0.25 69.1484063745022 ;
		END PORT
	END pin_65
	PIN pin_66
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 68.57868525896436 0.25 68.82868525896436 ;
		END PORT
	END pin_66
	PIN pin_67
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 68.25896414342651 0.25 68.50896414342651 ;
		END PORT
	END pin_67
	PIN pin_68
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 67.93924302788866 0.25 68.18924302788866 ;
		END PORT
	END pin_68
	PIN pin_69
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 67.61952191235082 0.25 67.86952191235082 ;
		END PORT
	END pin_69
	PIN pin_70
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 67.29980079681297 0.25 67.54980079681297 ;
		END PORT
	END pin_70
	PIN pin_71
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 66.98007968127513 0.25 67.23007968127513 ;
		END PORT
	END pin_71
	PIN pin_72
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 66.66035856573728 0.25 66.91035856573728 ;
		END PORT
	END pin_72
	PIN pin_73
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 66.34063745019944 0.25 66.59063745019944 ;
		END PORT
	END pin_73
	PIN pin_74
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 66.02091633466159 0.25 66.27091633466159 ;
		END PORT
	END pin_74
	PIN pin_75
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 65.70119521912375 0.25 65.95119521912375 ;
		END PORT
	END pin_75
	PIN pin_76
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 65.3814741035859 0.25 65.6314741035859 ;
		END PORT
	END pin_76
	PIN pin_77
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 65.06175298804806 0.25 65.31175298804806 ;
		END PORT
	END pin_77
	PIN pin_78
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 64.74203187251021 0.25 64.99203187251021 ;
		END PORT
	END pin_78
	PIN pin_79
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 64.42231075697237 0.25 64.67231075697237 ;
		END PORT
	END pin_79
	PIN pin_80
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 64.10258964143452 0.25 64.35258964143452 ;
		END PORT
	END pin_80
	PIN pin_81
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 63.782868525896674 0.25 64.03286852589667 ;
		END PORT
	END pin_81
	PIN pin_82
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 63.46314741035883 0.25 63.71314741035883 ;
		END PORT
	END pin_82
	PIN pin_83
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 63.14342629482098 0.25 63.39342629482098 ;
		END PORT
	END pin_83
	PIN pin_84
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 62.82370517928314 0.25 63.07370517928314 ;
		END PORT
	END pin_84
	PIN pin_85
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 62.50398406374529 0.25 62.75398406374529 ;
		END PORT
	END pin_85
	PIN pin_86
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 62.18426294820745 0.25 62.43426294820745 ;
		END PORT
	END pin_86
	PIN pin_87
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 61.8645418326696 0.25 62.1145418326696 ;
		END PORT
	END pin_87
	PIN pin_88
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 61.544820717131756 0.25 61.794820717131756 ;
		END PORT
	END pin_88
	PIN pin_89
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 61.22509960159391 0.25 61.47509960159391 ;
		END PORT
	END pin_89
	PIN pin_90
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 60.905378486056065 0.25 61.155378486056065 ;
		END PORT
	END pin_90
	PIN pin_91
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 60.58565737051822 0.25 60.83565737051822 ;
		END PORT
	END pin_91
	PIN pin_92
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 60.265936254980375 0.25 60.515936254980375 ;
		END PORT
	END pin_92
	PIN pin_93
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 59.94621513944253 0.25 60.19621513944253 ;
		END PORT
	END pin_93
	PIN pin_94
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 59.626494023904684 0.25 59.876494023904684 ;
		END PORT
	END pin_94
	PIN pin_95
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 59.30677290836684 0.25 59.55677290836684 ;
		END PORT
	END pin_95
	PIN pin_96
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.98705179282899 0.25 59.23705179282899 ;
		END PORT
	END pin_96
	PIN pin_97
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.66733067729115 0.25 58.91733067729115 ;
		END PORT
	END pin_97
	PIN pin_98
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.3476095617533 0.25 58.5976095617533 ;
		END PORT
	END pin_98
	PIN pin_99
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.02788844621546 0.25 58.27788844621546 ;
		END PORT
	END pin_99
	PIN pin_100
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 57.70816733067761 0.25 57.95816733067761 ;
		END PORT
	END pin_100
	PIN pin_101
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 57.388446215139766 0.25 57.638446215139766 ;
		END PORT
	END pin_101
	PIN pin_102
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 57.06872509960192 0.25 57.31872509960192 ;
		END PORT
	END pin_102
	PIN pin_103
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 56.749003984064075 0.25 56.999003984064075 ;
		END PORT
	END pin_103
	PIN pin_104
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 56.42928286852623 0.25 56.67928286852623 ;
		END PORT
	END pin_104
	PIN pin_105
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 56.109561752988384 0.25 56.359561752988384 ;
		END PORT
	END pin_105
	PIN pin_106
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 55.78984063745054 0.25 56.03984063745054 ;
		END PORT
	END pin_106
	PIN pin_107
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 55.47011952191269 0.25 55.72011952191269 ;
		END PORT
	END pin_107
	PIN pin_108
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 55.15039840637485 0.25 55.40039840637485 ;
		END PORT
	END pin_108
	PIN pin_109
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 54.830677290837 0.25 55.080677290837 ;
		END PORT
	END pin_109
	PIN pin_110
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 54.51095617529916 0.25 54.76095617529916 ;
		END PORT
	END pin_110
	PIN pin_111
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 54.19123505976131 0.25 54.44123505976131 ;
		END PORT
	END pin_111
	PIN pin_112
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 53.871513944223466 0.25 54.121513944223466 ;
		END PORT
	END pin_112
	PIN pin_113
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 53.55179282868562 0.25 53.80179282868562 ;
		END PORT
	END pin_113
	PIN pin_114
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 53.232071713147775 0.25 53.482071713147775 ;
		END PORT
	END pin_114
	PIN pin_115
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 52.91235059760993 0.25 53.16235059760993 ;
		END PORT
	END pin_115
	PIN pin_116
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 52.592629482072084 0.25 52.842629482072084 ;
		END PORT
	END pin_116
	PIN pin_117
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 52.27290836653424 0.25 52.52290836653424 ;
		END PORT
	END pin_117
	PIN pin_118
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 51.95318725099639 0.25 52.20318725099639 ;
		END PORT
	END pin_118
	PIN pin_119
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 51.63346613545855 0.25 51.88346613545855 ;
		END PORT
	END pin_119
	PIN pin_120
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 51.3137450199207 0.25 51.5637450199207 ;
		END PORT
	END pin_120
	PIN pin_121
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 50.99402390438286 0.25 51.24402390438286 ;
		END PORT
	END pin_121
	PIN pin_122
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 50.67430278884501 0.25 50.92430278884501 ;
		END PORT
	END pin_122
	PIN pin_123
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 50.354581673307166 0.25 50.604581673307166 ;
		END PORT
	END pin_123
	PIN pin_124
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 50.03486055776932 0.25 50.28486055776932 ;
		END PORT
	END pin_124
	PIN pin_125
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 49.715139442231475 0.25 49.965139442231475 ;
		END PORT
	END pin_125
	PIN pin_126
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 49.39541832669363 0.25 49.64541832669363 ;
		END PORT
	END pin_126
	PIN pin_127
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 49.075697211155784 0.25 49.325697211155784 ;
		END PORT
	END pin_127
	PIN pin_128
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 48.75597609561794 0.25 49.00597609561794 ;
		END PORT
	END pin_128
	PIN pin_129
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 48.43625498008009 0.25 48.68625498008009 ;
		END PORT
	END pin_129
	PIN pin_130
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 48.11653386454225 0.25 48.36653386454225 ;
		END PORT
	END pin_130
	PIN pin_131
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 47.7968127490044 0.25 48.0468127490044 ;
		END PORT
	END pin_131
	PIN pin_132
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 47.47709163346656 0.25 47.72709163346656 ;
		END PORT
	END pin_132
	PIN pin_133
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 47.15737051792871 0.25 47.40737051792871 ;
		END PORT
	END pin_133
	PIN pin_134
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 46.837649402390866 0.25 47.087649402390866 ;
		END PORT
	END pin_134
	PIN pin_135
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 46.51792828685302 0.25 46.76792828685302 ;
		END PORT
	END pin_135
	PIN pin_136
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 46.198207171315175 0.25 46.448207171315175 ;
		END PORT
	END pin_136
	PIN pin_137
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 45.87848605577733 0.25 46.12848605577733 ;
		END PORT
	END pin_137
	PIN pin_138
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 45.558764940239485 0.25 45.808764940239485 ;
		END PORT
	END pin_138
	PIN pin_139
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 45.23904382470164 0.25 45.48904382470164 ;
		END PORT
	END pin_139
	PIN pin_140
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 44.919322709163794 0.25 45.169322709163794 ;
		END PORT
	END pin_140
	PIN pin_141
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 44.59960159362595 0.25 44.84960159362595 ;
		END PORT
	END pin_141
	PIN pin_142
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 44.2798804780881 0.25 44.5298804780881 ;
		END PORT
	END pin_142
	PIN pin_143
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 43.96015936255026 0.25 44.21015936255026 ;
		END PORT
	END pin_143
	PIN pin_144
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 43.64043824701241 0.25 43.89043824701241 ;
		END PORT
	END pin_144
	PIN pin_145
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 43.32071713147457 0.25 43.57071713147457 ;
		END PORT
	END pin_145
	PIN pin_146
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 43.00099601593672 0.25 43.25099601593672 ;
		END PORT
	END pin_146
	PIN pin_147
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 42.681274900398876 0.25 42.931274900398876 ;
		END PORT
	END pin_147
	PIN pin_148
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 42.36155378486103 0.25 42.61155378486103 ;
		END PORT
	END pin_148
	PIN pin_149
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 42.041832669323185 0.25 42.291832669323185 ;
		END PORT
	END pin_149
	PIN pin_150
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 41.72211155378534 0.25 41.97211155378534 ;
		END PORT
	END pin_150
	PIN pin_151
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 41.402390438247494 0.25 41.652390438247494 ;
		END PORT
	END pin_151
	PIN pin_152
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 41.08266932270965 0.25 41.33266932270965 ;
		END PORT
	END pin_152
	PIN pin_153
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 40.7629482071718 0.25 41.0129482071718 ;
		END PORT
	END pin_153
	PIN pin_154
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 40.44322709163396 0.25 40.69322709163396 ;
		END PORT
	END pin_154
	PIN pin_155
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 40.12350597609611 0.25 40.37350597609611 ;
		END PORT
	END pin_155
	PIN pin_156
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 39.80378486055827 0.25 40.05378486055827 ;
		END PORT
	END pin_156
	PIN pin_157
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 39.48406374502042 0.25 39.73406374502042 ;
		END PORT
	END pin_157
	PIN pin_158
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 39.164342629482576 0.25 39.414342629482576 ;
		END PORT
	END pin_158
	PIN pin_159
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 38.84462151394473 0.25 39.09462151394473 ;
		END PORT
	END pin_159
	PIN pin_160
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 38.524900398406885 0.25 38.774900398406885 ;
		END PORT
	END pin_160
	PIN pin_161
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 38.20517928286904 0.25 38.45517928286904 ;
		END PORT
	END pin_161
	PIN pin_162
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 37.885458167331194 0.25 38.135458167331194 ;
		END PORT
	END pin_162
	PIN pin_163
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 37.56573705179335 0.25 37.81573705179335 ;
		END PORT
	END pin_163
	PIN pin_164
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 37.2460159362555 0.25 37.4960159362555 ;
		END PORT
	END pin_164
	PIN pin_165
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 36.92629482071766 0.25 37.17629482071766 ;
		END PORT
	END pin_165
	PIN pin_166
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 36.60657370517981 0.25 36.85657370517981 ;
		END PORT
	END pin_166
	PIN pin_167
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 36.28685258964197 0.25 36.53685258964197 ;
		END PORT
	END pin_167
	PIN pin_168
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 35.96713147410412 0.25 36.21713147410412 ;
		END PORT
	END pin_168
	PIN pin_169
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 35.647410358566276 0.25 35.897410358566276 ;
		END PORT
	END pin_169
	PIN pin_170
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 35.32768924302843 0.25 35.57768924302843 ;
		END PORT
	END pin_170
	PIN pin_171
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 35.007968127490585 0.25 35.257968127490585 ;
		END PORT
	END pin_171
	PIN pin_172
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 34.68824701195274 0.25 34.93824701195274 ;
		END PORT
	END pin_172
	PIN pin_173
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 34.368525896414894 0.25 34.618525896414894 ;
		END PORT
	END pin_173
	PIN pin_174
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 34.04880478087705 0.25 34.29880478087705 ;
		END PORT
	END pin_174
	PIN pin_175
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 33.7290836653392 0.25 33.9790836653392 ;
		END PORT
	END pin_175
	PIN pin_176
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 33.40936254980136 0.25 33.65936254980136 ;
		END PORT
	END pin_176
	PIN pin_177
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 33.08964143426351 0.25 33.33964143426351 ;
		END PORT
	END pin_177
	PIN pin_178
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 32.76992031872567 0.25 33.01992031872567 ;
		END PORT
	END pin_178
	PIN pin_179
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 32.45019920318782 0.25 32.70019920318782 ;
		END PORT
	END pin_179
	PIN pin_180
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 32.130478087649976 0.25 32.380478087649976 ;
		END PORT
	END pin_180
	PIN pin_181
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 31.81075697211213 0.25 32.06075697211213 ;
		END PORT
	END pin_181
	PIN pin_182
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 31.491035856574282 0.25 31.741035856574282 ;
		END PORT
	END pin_182
	PIN pin_183
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 31.171314741036433 0.25 31.421314741036433 ;
		END PORT
	END pin_183
	PIN pin_184
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 30.851593625498584 0.25 31.101593625498584 ;
		END PORT
	END pin_184
	PIN pin_185
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 30.531872509960735 0.25 30.781872509960735 ;
		END PORT
	END pin_185
	PIN pin_186
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 30.212151394422886 0.25 30.462151394422886 ;
		END PORT
	END pin_186
	PIN pin_187
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 29.892430278885037 0.25 30.142430278885037 ;
		END PORT
	END pin_187
	PIN pin_188
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 29.572709163347188 0.25 29.822709163347188 ;
		END PORT
	END pin_188
	PIN pin_189
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 29.25298804780934 0.25 29.50298804780934 ;
		END PORT
	END pin_189
	PIN pin_190
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 28.93326693227149 0.25 29.18326693227149 ;
		END PORT
	END pin_190
	PIN pin_191
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 28.61354581673364 0.25 28.86354581673364 ;
		END PORT
	END pin_191
	PIN pin_192
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 28.293824701195792 0.25 28.543824701195792 ;
		END PORT
	END pin_192
	PIN pin_193
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 27.974103585657943 0.25 28.224103585657943 ;
		END PORT
	END pin_193
	PIN pin_194
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 27.654382470120094 0.25 27.904382470120094 ;
		END PORT
	END pin_194
	PIN pin_195
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 27.334661354582245 0.25 27.584661354582245 ;
		END PORT
	END pin_195
	PIN pin_196
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 27.014940239044396 0.25 27.264940239044396 ;
		END PORT
	END pin_196
	PIN pin_197
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 26.695219123506547 0.25 26.945219123506547 ;
		END PORT
	END pin_197
	PIN pin_198
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 26.375498007968698 0.25 26.625498007968698 ;
		END PORT
	END pin_198
	PIN pin_199
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 26.05577689243085 0.25 26.30577689243085 ;
		END PORT
	END pin_199
	PIN pin_200
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 25.736055776893 0.25 25.986055776893 ;
		END PORT
	END pin_200
	PIN pin_201
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 25.41633466135515 0.25 25.66633466135515 ;
		END PORT
	END pin_201
	PIN pin_202
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 25.096613545817302 0.25 25.346613545817302 ;
		END PORT
	END pin_202
	PIN pin_203
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 24.776892430279453 0.25 25.026892430279453 ;
		END PORT
	END pin_203
	PIN pin_204
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 24.457171314741604 0.25 24.707171314741604 ;
		END PORT
	END pin_204
	PIN pin_205
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 24.137450199203755 0.25 24.387450199203755 ;
		END PORT
	END pin_205
	PIN pin_206
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 23.817729083665906 0.25 24.067729083665906 ;
		END PORT
	END pin_206
	PIN pin_207
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 23.498007968128057 0.25 23.748007968128057 ;
		END PORT
	END pin_207
	PIN pin_208
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 23.178286852590208 0.25 23.428286852590208 ;
		END PORT
	END pin_208
	PIN pin_209
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 22.85856573705236 0.25 23.10856573705236 ;
		END PORT
	END pin_209
	PIN pin_210
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 22.53884462151451 0.25 22.78884462151451 ;
		END PORT
	END pin_210
	PIN pin_211
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 22.21912350597666 0.25 22.46912350597666 ;
		END PORT
	END pin_211
	PIN pin_212
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 21.899402390438812 0.25 22.149402390438812 ;
		END PORT
	END pin_212
	PIN pin_213
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 21.579681274900963 0.25 21.829681274900963 ;
		END PORT
	END pin_213
	PIN pin_214
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 21.259960159363114 0.25 21.509960159363114 ;
		END PORT
	END pin_214
	PIN pin_215
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 20.940239043825265 0.25 21.190239043825265 ;
		END PORT
	END pin_215
	PIN pin_216
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 20.620517928287416 0.25 20.870517928287416 ;
		END PORT
	END pin_216
	PIN pin_217
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 20.300796812749567 0.25 20.550796812749567 ;
		END PORT
	END pin_217
	PIN pin_218
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 19.98107569721172 0.25 20.23107569721172 ;
		END PORT
	END pin_218
	PIN pin_219
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 19.66135458167387 0.25 19.91135458167387 ;
		END PORT
	END pin_219
	PIN pin_220
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 19.34163346613602 0.25 19.59163346613602 ;
		END PORT
	END pin_220
	PIN pin_221
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 19.02191235059817 0.25 19.27191235059817 ;
		END PORT
	END pin_221
	PIN pin_222
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 18.702191235060322 0.25 18.952191235060322 ;
		END PORT
	END pin_222
	PIN pin_223
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 18.382470119522473 0.25 18.632470119522473 ;
		END PORT
	END pin_223
	PIN pin_224
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 18.062749003984624 0.25 18.312749003984624 ;
		END PORT
	END pin_224
	PIN pin_225
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 17.743027888446775 0.25 17.993027888446775 ;
		END PORT
	END pin_225
	PIN pin_226
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 17.423306772908926 0.25 17.673306772908926 ;
		END PORT
	END pin_226
	PIN pin_227
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 17.103585657371077 0.25 17.353585657371077 ;
		END PORT
	END pin_227
	PIN pin_228
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 16.78386454183323 0.25 17.03386454183323 ;
		END PORT
	END pin_228
	PIN pin_229
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 16.46414342629538 0.25 16.71414342629538 ;
		END PORT
	END pin_229
	PIN pin_230
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 16.14442231075753 0.25 16.39442231075753 ;
		END PORT
	END pin_230
	PIN pin_231
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 15.824701195219681 0.25 16.07470119521968 ;
		END PORT
	END pin_231
	PIN pin_232
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 15.504980079681832 0.25 15.754980079681832 ;
		END PORT
	END pin_232
	PIN pin_233
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 15.185258964143983 0.25 15.435258964143983 ;
		END PORT
	END pin_233
	PIN pin_234
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 14.865537848606134 0.25 15.115537848606134 ;
		END PORT
	END pin_234
	PIN pin_235
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 14.545816733068285 0.25 14.795816733068285 ;
		END PORT
	END pin_235
	PIN pin_236
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 14.226095617530436 0.25 14.476095617530436 ;
		END PORT
	END pin_236
	PIN pin_237
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 13.906374501992588 0.25 14.156374501992588 ;
		END PORT
	END pin_237
	PIN pin_238
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 13.586653386454739 0.25 13.836653386454739 ;
		END PORT
	END pin_238
	PIN pin_239
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 13.26693227091689 0.25 13.51693227091689 ;
		END PORT
	END pin_239
	PIN pin_240
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 12.94721115537904 0.25 13.19721115537904 ;
		END PORT
	END pin_240
	PIN pin_241
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 12.627490039841192 0.25 12.877490039841192 ;
		END PORT
	END pin_241
	PIN pin_242
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 12.307768924303343 0.25 12.557768924303343 ;
		END PORT
	END pin_242
	PIN pin_243
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 11.988047808765494 0.25 12.238047808765494 ;
		END PORT
	END pin_243
	PIN pin_244
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 11.668326693227645 0.25 11.918326693227645 ;
		END PORT
	END pin_244
	PIN pin_245
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 11.348605577689796 0.25 11.598605577689796 ;
		END PORT
	END pin_245
	PIN pin_246
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 11.028884462151947 0.25 11.278884462151947 ;
		END PORT
	END pin_246
	PIN pin_247
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 10.709163346614098 0.25 10.959163346614098 ;
		END PORT
	END pin_247
	PIN pin_248
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 10.389442231076249 0.25 10.639442231076249 ;
		END PORT
	END pin_248
	PIN pin_249
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 10.0697211155384 0.25 10.3197211155384 ;
		END PORT
	END pin_249
	PIN pin_250
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.069721115537849 100 10.319721115537849 ;
		END PORT
	END pin_250
	PIN pin_251
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.389442231075698 100 10.639442231075698 ;
		END PORT
	END pin_251
	PIN pin_252
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.709163346613547 100 10.959163346613547 ;
		END PORT
	END pin_252
	PIN pin_253
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.028884462151396 100 11.278884462151396 ;
		END PORT
	END pin_253
	PIN pin_254
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.348605577689245 100 11.598605577689245 ;
		END PORT
	END pin_254
	PIN pin_255
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.668326693227094 100 11.918326693227094 ;
		END PORT
	END pin_255
	PIN pin_256
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.988047808764943 100 12.238047808764943 ;
		END PORT
	END pin_256
	PIN pin_257
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.307768924302792 100 12.557768924302792 ;
		END PORT
	END pin_257
	PIN pin_258
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.627490039840641 100 12.877490039840641 ;
		END PORT
	END pin_258
	PIN pin_259
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.94721115537849 100 13.19721115537849 ;
		END PORT
	END pin_259
	PIN pin_260
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.266932270916339 100 13.516932270916339 ;
		END PORT
	END pin_260
	PIN pin_261
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.586653386454188 100 13.836653386454188 ;
		END PORT
	END pin_261
	PIN pin_262
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.906374501992037 100 14.156374501992037 ;
		END PORT
	END pin_262
	PIN pin_263
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.226095617529886 100 14.476095617529886 ;
		END PORT
	END pin_263
	PIN pin_264
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.545816733067735 100 14.795816733067735 ;
		END PORT
	END pin_264
	PIN pin_265
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.865537848605584 100 15.115537848605584 ;
		END PORT
	END pin_265
	PIN pin_266
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.185258964143433 100 15.435258964143433 ;
		END PORT
	END pin_266
	PIN pin_267
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.504980079681282 100 15.754980079681282 ;
		END PORT
	END pin_267
	PIN pin_268
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.82470119521913 100 16.07470119521913 ;
		END PORT
	END pin_268
	PIN pin_269
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.14442231075698 100 16.39442231075698 ;
		END PORT
	END pin_269
	PIN pin_270
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.46414342629483 100 16.71414342629483 ;
		END PORT
	END pin_270
	PIN pin_271
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.783864541832678 100 17.033864541832678 ;
		END PORT
	END pin_271
	PIN pin_272
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.103585657370527 100 17.353585657370527 ;
		END PORT
	END pin_272
	PIN pin_273
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.423306772908376 100 17.673306772908376 ;
		END PORT
	END pin_273
	PIN pin_274
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.743027888446225 100 17.993027888446225 ;
		END PORT
	END pin_274
	PIN pin_275
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.062749003984074 100 18.312749003984074 ;
		END PORT
	END pin_275
	PIN pin_276
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.382470119521923 100 18.632470119521923 ;
		END PORT
	END pin_276
	PIN pin_277
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.70219123505977 100 18.95219123505977 ;
		END PORT
	END pin_277
	PIN pin_278
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.02191235059762 100 19.27191235059762 ;
		END PORT
	END pin_278
	PIN pin_279
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.34163346613547 100 19.59163346613547 ;
		END PORT
	END pin_279
	PIN pin_280
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.66135458167332 100 19.91135458167332 ;
		END PORT
	END pin_280
	PIN pin_281
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.981075697211168 100 20.231075697211168 ;
		END PORT
	END pin_281
	PIN pin_282
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.300796812749017 100 20.550796812749017 ;
		END PORT
	END pin_282
	PIN pin_283
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.620517928286866 100 20.870517928286866 ;
		END PORT
	END pin_283
	PIN pin_284
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.940239043824715 100 21.190239043824715 ;
		END PORT
	END pin_284
	PIN pin_285
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.259960159362564 100 21.509960159362564 ;
		END PORT
	END pin_285
	PIN pin_286
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.579681274900413 100 21.829681274900413 ;
		END PORT
	END pin_286
	PIN pin_287
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.89940239043826 100 22.14940239043826 ;
		END PORT
	END pin_287
	PIN pin_288
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.21912350597611 100 22.46912350597611 ;
		END PORT
	END pin_288
	PIN pin_289
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.53884462151396 100 22.78884462151396 ;
		END PORT
	END pin_289
	PIN pin_290
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.85856573705181 100 23.10856573705181 ;
		END PORT
	END pin_290
	PIN pin_291
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.178286852589657 100 23.428286852589657 ;
		END PORT
	END pin_291
	PIN pin_292
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.498007968127506 100 23.748007968127506 ;
		END PORT
	END pin_292
	PIN pin_293
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.817729083665355 100 24.067729083665355 ;
		END PORT
	END pin_293
	PIN pin_294
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.137450199203204 100 24.387450199203204 ;
		END PORT
	END pin_294
	PIN pin_295
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.457171314741053 100 24.707171314741053 ;
		END PORT
	END pin_295
	PIN pin_296
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.776892430278902 100 25.026892430278902 ;
		END PORT
	END pin_296
	PIN pin_297
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.09661354581675 100 25.34661354581675 ;
		END PORT
	END pin_297
	PIN pin_298
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.4163346613546 100 25.6663346613546 ;
		END PORT
	END pin_298
	PIN pin_299
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.73605577689245 100 25.98605577689245 ;
		END PORT
	END pin_299
	PIN pin_300
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.0557768924303 100 26.3057768924303 ;
		END PORT
	END pin_300
	PIN pin_301
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.375498007968147 100 26.625498007968147 ;
		END PORT
	END pin_301
	PIN pin_302
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.695219123505996 100 26.945219123505996 ;
		END PORT
	END pin_302
	PIN pin_303
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.014940239043845 100 27.264940239043845 ;
		END PORT
	END pin_303
	PIN pin_304
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.334661354581694 100 27.584661354581694 ;
		END PORT
	END pin_304
	PIN pin_305
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.654382470119543 100 27.904382470119543 ;
		END PORT
	END pin_305
	PIN pin_306
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.974103585657392 100 28.224103585657392 ;
		END PORT
	END pin_306
	PIN pin_307
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.29382470119524 100 28.54382470119524 ;
		END PORT
	END pin_307
	PIN pin_308
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.61354581673309 100 28.86354581673309 ;
		END PORT
	END pin_308
	PIN pin_309
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.93326693227094 100 29.18326693227094 ;
		END PORT
	END pin_309
	PIN pin_310
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.25298804780879 100 29.50298804780879 ;
		END PORT
	END pin_310
	PIN pin_311
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.572709163346637 100 29.822709163346637 ;
		END PORT
	END pin_311
	PIN pin_312
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.892430278884486 100 30.142430278884486 ;
		END PORT
	END pin_312
	PIN pin_313
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.212151394422335 100 30.462151394422335 ;
		END PORT
	END pin_313
	PIN pin_314
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.531872509960184 100 30.781872509960184 ;
		END PORT
	END pin_314
	PIN pin_315
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.851593625498033 100 31.101593625498033 ;
		END PORT
	END pin_315
	PIN pin_316
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.171314741035882 100 31.421314741035882 ;
		END PORT
	END pin_316
	PIN pin_317
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.49103585657373 100 31.74103585657373 ;
		END PORT
	END pin_317
	PIN pin_318
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.81075697211158 100 32.06075697211158 ;
		END PORT
	END pin_318
	PIN pin_319
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.13047808764942 100 32.38047808764942 ;
		END PORT
	END pin_319
	PIN pin_320
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.45019920318727 100 32.70019920318727 ;
		END PORT
	END pin_320
	PIN pin_321
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.76992031872511 100 33.01992031872511 ;
		END PORT
	END pin_321
	PIN pin_322
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.08964143426296 100 33.33964143426296 ;
		END PORT
	END pin_322
	PIN pin_323
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.409362549800804 100 33.659362549800804 ;
		END PORT
	END pin_323
	PIN pin_324
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.72908366533865 100 33.97908366533865 ;
		END PORT
	END pin_324
	PIN pin_325
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.048804780876495 100 34.298804780876495 ;
		END PORT
	END pin_325
	PIN pin_326
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.36852589641434 100 34.61852589641434 ;
		END PORT
	END pin_326
	PIN pin_327
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.688247011952186 100 34.938247011952186 ;
		END PORT
	END pin_327
	PIN pin_328
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.00796812749003 100 35.25796812749003 ;
		END PORT
	END pin_328
	PIN pin_329
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.327689243027876 100 35.577689243027876 ;
		END PORT
	END pin_329
	PIN pin_330
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.64741035856572 100 35.89741035856572 ;
		END PORT
	END pin_330
	PIN pin_331
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.96713147410357 100 36.21713147410357 ;
		END PORT
	END pin_331
	PIN pin_332
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.28685258964141 100 36.53685258964141 ;
		END PORT
	END pin_332
	PIN pin_333
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.60657370517926 100 36.85657370517926 ;
		END PORT
	END pin_333
	PIN pin_334
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.926294820717104 100 37.176294820717104 ;
		END PORT
	END pin_334
	PIN pin_335
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.24601593625495 100 37.49601593625495 ;
		END PORT
	END pin_335
	PIN pin_336
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.565737051792794 100 37.815737051792794 ;
		END PORT
	END pin_336
	PIN pin_337
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.88545816733064 100 38.13545816733064 ;
		END PORT
	END pin_337
	PIN pin_338
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.205179282868485 100 38.455179282868485 ;
		END PORT
	END pin_338
	PIN pin_339
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.52490039840633 100 38.77490039840633 ;
		END PORT
	END pin_339
	PIN pin_340
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.844621513944176 100 39.094621513944176 ;
		END PORT
	END pin_340
	PIN pin_341
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.16434262948202 100 39.41434262948202 ;
		END PORT
	END pin_341
	PIN pin_342
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.48406374501987 100 39.73406374501987 ;
		END PORT
	END pin_342
	PIN pin_343
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.80378486055771 100 40.05378486055771 ;
		END PORT
	END pin_343
	PIN pin_344
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.12350597609556 100 40.37350597609556 ;
		END PORT
	END pin_344
	PIN pin_345
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.4432270916334 100 40.6932270916334 ;
		END PORT
	END pin_345
	PIN pin_346
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.76294820717125 100 41.01294820717125 ;
		END PORT
	END pin_346
	PIN pin_347
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.082669322709094 100 41.332669322709094 ;
		END PORT
	END pin_347
	PIN pin_348
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.40239043824694 100 41.65239043824694 ;
		END PORT
	END pin_348
	PIN pin_349
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.722111553784785 100 41.972111553784785 ;
		END PORT
	END pin_349
	PIN pin_350
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.04183266932263 100 42.29183266932263 ;
		END PORT
	END pin_350
	PIN pin_351
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.361553784860476 100 42.611553784860476 ;
		END PORT
	END pin_351
	PIN pin_352
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.68127490039832 100 42.93127490039832 ;
		END PORT
	END pin_352
	PIN pin_353
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.00099601593617 100 43.25099601593617 ;
		END PORT
	END pin_353
	PIN pin_354
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.32071713147401 100 43.57071713147401 ;
		END PORT
	END pin_354
	PIN pin_355
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.64043824701186 100 43.89043824701186 ;
		END PORT
	END pin_355
	PIN pin_356
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.9601593625497 100 44.2101593625497 ;
		END PORT
	END pin_356
	PIN pin_357
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.27988047808755 100 44.52988047808755 ;
		END PORT
	END pin_357
	PIN pin_358
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.599601593625394 100 44.849601593625394 ;
		END PORT
	END pin_358
	PIN pin_359
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.91932270916324 100 45.16932270916324 ;
		END PORT
	END pin_359
	PIN pin_360
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.239043824701085 100 45.489043824701085 ;
		END PORT
	END pin_360
	PIN pin_361
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.55876494023893 100 45.80876494023893 ;
		END PORT
	END pin_361
	PIN pin_362
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.878486055776776 100 46.128486055776776 ;
		END PORT
	END pin_362
	PIN pin_363
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.19820717131462 100 46.44820717131462 ;
		END PORT
	END pin_363
	PIN pin_364
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.51792828685247 100 46.76792828685247 ;
		END PORT
	END pin_364
	PIN pin_365
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.83764940239031 100 47.08764940239031 ;
		END PORT
	END pin_365
	PIN pin_366
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.15737051792816 100 47.40737051792816 ;
		END PORT
	END pin_366
	PIN pin_367
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.477091633466 100 47.727091633466 ;
		END PORT
	END pin_367
	PIN pin_368
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.79681274900385 100 48.04681274900385 ;
		END PORT
	END pin_368
	PIN pin_369
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.116533864541694 100 48.366533864541694 ;
		END PORT
	END pin_369
	PIN pin_370
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.43625498007954 100 48.68625498007954 ;
		END PORT
	END pin_370
	PIN pin_371
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.755976095617385 100 49.005976095617385 ;
		END PORT
	END pin_371
	PIN pin_372
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.07569721115523 100 49.32569721115523 ;
		END PORT
	END pin_372
	PIN pin_373
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.395418326693076 100 49.645418326693076 ;
		END PORT
	END pin_373
	PIN pin_374
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.71513944223092 100 49.96513944223092 ;
		END PORT
	END pin_374
	PIN pin_375
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.034860557768766 100 50.284860557768766 ;
		END PORT
	END pin_375
	PIN pin_376
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.35458167330661 100 50.60458167330661 ;
		END PORT
	END pin_376
	PIN pin_377
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.67430278884446 100 50.92430278884446 ;
		END PORT
	END pin_377
	PIN pin_378
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.9940239043823 100 51.2440239043823 ;
		END PORT
	END pin_378
	PIN pin_379
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.31374501992015 100 51.56374501992015 ;
		END PORT
	END pin_379
	PIN pin_380
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.633466135457994 100 51.883466135457994 ;
		END PORT
	END pin_380
	PIN pin_381
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.95318725099584 100 52.20318725099584 ;
		END PORT
	END pin_381
	PIN pin_382
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.272908366533684 100 52.522908366533684 ;
		END PORT
	END pin_382
	PIN pin_383
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.59262948207153 100 52.84262948207153 ;
		END PORT
	END pin_383
	PIN pin_384
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.912350597609375 100 53.162350597609375 ;
		END PORT
	END pin_384
	PIN pin_385
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.23207171314722 100 53.48207171314722 ;
		END PORT
	END pin_385
	PIN pin_386
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.551792828685066 100 53.801792828685066 ;
		END PORT
	END pin_386
	PIN pin_387
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.87151394422291 100 54.12151394422291 ;
		END PORT
	END pin_387
	PIN pin_388
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.19123505976076 100 54.44123505976076 ;
		END PORT
	END pin_388
	PIN pin_389
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.5109561752986 100 54.7609561752986 ;
		END PORT
	END pin_389
	PIN pin_390
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.83067729083645 100 55.08067729083645 ;
		END PORT
	END pin_390
	PIN pin_391
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.15039840637429 100 55.40039840637429 ;
		END PORT
	END pin_391
	PIN pin_392
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.47011952191214 100 55.72011952191214 ;
		END PORT
	END pin_392
	PIN pin_393
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.789840637449984 100 56.039840637449984 ;
		END PORT
	END pin_393
	PIN pin_394
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.10956175298783 100 56.35956175298783 ;
		END PORT
	END pin_394
	PIN pin_395
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.429282868525675 100 56.679282868525675 ;
		END PORT
	END pin_395
	PIN pin_396
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.74900398406352 100 56.99900398406352 ;
		END PORT
	END pin_396
	PIN pin_397
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.068725099601366 100 57.318725099601366 ;
		END PORT
	END pin_397
	PIN pin_398
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.38844621513921 100 57.63844621513921 ;
		END PORT
	END pin_398
	PIN pin_399
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.70816733067706 100 57.95816733067706 ;
		END PORT
	END pin_399
	PIN pin_400
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.0278884462149 100 58.2778884462149 ;
		END PORT
	END pin_400
	PIN pin_401
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.34760956175275 100 58.59760956175275 ;
		END PORT
	END pin_401
	PIN pin_402
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.66733067729059 100 58.91733067729059 ;
		END PORT
	END pin_402
	PIN pin_403
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.98705179282844 100 59.23705179282844 ;
		END PORT
	END pin_403
	PIN pin_404
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.306772908366284 100 59.556772908366284 ;
		END PORT
	END pin_404
	PIN pin_405
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.62649402390413 100 59.87649402390413 ;
		END PORT
	END pin_405
	PIN pin_406
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.946215139441975 100 60.196215139441975 ;
		END PORT
	END pin_406
	PIN pin_407
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.26593625497982 100 60.51593625497982 ;
		END PORT
	END pin_407
	PIN pin_408
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.585657370517666 100 60.835657370517666 ;
		END PORT
	END pin_408
	PIN pin_409
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.90537848605551 100 61.15537848605551 ;
		END PORT
	END pin_409
	PIN pin_410
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.22509960159336 100 61.47509960159336 ;
		END PORT
	END pin_410
	PIN pin_411
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.5448207171312 100 61.7948207171312 ;
		END PORT
	END pin_411
	PIN pin_412
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.86454183266905 100 62.11454183266905 ;
		END PORT
	END pin_412
	PIN pin_413
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.18426294820689 100 62.43426294820689 ;
		END PORT
	END pin_413
	PIN pin_414
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.50398406374474 100 62.75398406374474 ;
		END PORT
	END pin_414
	PIN pin_415
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.823705179282584 100 63.073705179282584 ;
		END PORT
	END pin_415
	PIN pin_416
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.14342629482043 100 63.39342629482043 ;
		END PORT
	END pin_416
	PIN pin_417
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.463147410358275 100 63.713147410358275 ;
		END PORT
	END pin_417
	PIN pin_418
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.78286852589612 100 64.03286852589612 ;
		END PORT
	END pin_418
	PIN pin_419
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.10258964143397 100 64.35258964143397 ;
		END PORT
	END pin_419
	PIN pin_420
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.42231075697181 100 64.67231075697181 ;
		END PORT
	END pin_420
	PIN pin_421
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.74203187250966 100 64.99203187250966 ;
		END PORT
	END pin_421
	PIN pin_422
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.0617529880475 100 65.3117529880475 ;
		END PORT
	END pin_422
	PIN pin_423
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.38147410358535 100 65.63147410358535 ;
		END PORT
	END pin_423
	PIN pin_424
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.70119521912319 100 65.95119521912319 ;
		END PORT
	END pin_424
	PIN pin_425
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.02091633466104 100 66.27091633466104 ;
		END PORT
	END pin_425
	PIN pin_426
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.34063745019888 100 66.59063745019888 ;
		END PORT
	END pin_426
	PIN pin_427
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.66035856573673 100 66.91035856573673 ;
		END PORT
	END pin_427
	PIN pin_428
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.98007968127457 100 67.23007968127457 ;
		END PORT
	END pin_428
	PIN pin_429
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.29980079681242 100 67.54980079681242 ;
		END PORT
	END pin_429
	PIN pin_430
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.61952191235027 100 67.86952191235027 ;
		END PORT
	END pin_430
	PIN pin_431
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.93924302788811 100 68.18924302788811 ;
		END PORT
	END pin_431
	PIN pin_432
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.25896414342596 100 68.50896414342596 ;
		END PORT
	END pin_432
	PIN pin_433
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.5786852589638 100 68.8286852589638 ;
		END PORT
	END pin_433
	PIN pin_434
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.89840637450165 100 69.14840637450165 ;
		END PORT
	END pin_434
	PIN pin_435
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.21812749003949 100 69.46812749003949 ;
		END PORT
	END pin_435
	PIN pin_436
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.53784860557734 100 69.78784860557734 ;
		END PORT
	END pin_436
	PIN pin_437
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.85756972111518 100 70.10756972111518 ;
		END PORT
	END pin_437
	PIN pin_438
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.17729083665303 100 70.42729083665303 ;
		END PORT
	END pin_438
	PIN pin_439
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.49701195219087 100 70.74701195219087 ;
		END PORT
	END pin_439
	PIN pin_440
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.81673306772872 100 71.06673306772872 ;
		END PORT
	END pin_440
	PIN pin_441
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.13645418326657 100 71.38645418326657 ;
		END PORT
	END pin_441
	PIN pin_442
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.45617529880441 100 71.70617529880441 ;
		END PORT
	END pin_442
	PIN pin_443
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.77589641434226 100 72.02589641434226 ;
		END PORT
	END pin_443
	PIN pin_444
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.0956175298801 100 72.3456175298801 ;
		END PORT
	END pin_444
	PIN pin_445
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.41533864541795 100 72.66533864541795 ;
		END PORT
	END pin_445
	PIN pin_446
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.73505976095579 100 72.98505976095579 ;
		END PORT
	END pin_446
	PIN pin_447
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.05478087649364 100 73.30478087649364 ;
		END PORT
	END pin_447
	PIN pin_448
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.37450199203148 100 73.62450199203148 ;
		END PORT
	END pin_448
	PIN pin_449
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.69422310756933 100 73.94422310756933 ;
		END PORT
	END pin_449
	PIN pin_450
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.01394422310717 100 74.26394422310717 ;
		END PORT
	END pin_450
	PIN pin_451
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.33366533864502 100 74.58366533864502 ;
		END PORT
	END pin_451
	PIN pin_452
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.65338645418286 100 74.90338645418286 ;
		END PORT
	END pin_452
	PIN pin_453
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.97310756972071 100 75.22310756972071 ;
		END PORT
	END pin_453
	PIN pin_454
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.29282868525856 100 75.54282868525856 ;
		END PORT
	END pin_454
	PIN pin_455
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.6125498007964 100 75.8625498007964 ;
		END PORT
	END pin_455
	PIN pin_456
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.93227091633425 100 76.18227091633425 ;
		END PORT
	END pin_456
	PIN pin_457
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.25199203187209 100 76.50199203187209 ;
		END PORT
	END pin_457
	PIN pin_458
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.57171314740994 100 76.82171314740994 ;
		END PORT
	END pin_458
	PIN pin_459
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.89143426294778 100 77.14143426294778 ;
		END PORT
	END pin_459
	PIN pin_460
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.21115537848563 100 77.46115537848563 ;
		END PORT
	END pin_460
	PIN pin_461
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.53087649402347 100 77.78087649402347 ;
		END PORT
	END pin_461
	PIN pin_462
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.85059760956132 100 78.10059760956132 ;
		END PORT
	END pin_462
	PIN pin_463
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.17031872509916 100 78.42031872509916 ;
		END PORT
	END pin_463
	PIN pin_464
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.49003984063701 100 78.74003984063701 ;
		END PORT
	END pin_464
	PIN pin_465
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.80976095617486 100 79.05976095617486 ;
		END PORT
	END pin_465
	PIN pin_466
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.1294820717127 100 79.3794820717127 ;
		END PORT
	END pin_466
	PIN pin_467
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.44920318725055 100 79.69920318725055 ;
		END PORT
	END pin_467
	PIN pin_468
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.76892430278839 100 80.01892430278839 ;
		END PORT
	END pin_468
	PIN pin_469
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.08864541832624 100 80.33864541832624 ;
		END PORT
	END pin_469
	PIN pin_470
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.40836653386408 100 80.65836653386408 ;
		END PORT
	END pin_470
	PIN pin_471
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.72808764940193 100 80.97808764940193 ;
		END PORT
	END pin_471
	PIN pin_472
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.04780876493977 100 81.29780876493977 ;
		END PORT
	END pin_472
	PIN pin_473
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.36752988047762 100 81.61752988047762 ;
		END PORT
	END pin_473
	PIN pin_474
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.68725099601546 100 81.93725099601546 ;
		END PORT
	END pin_474
	PIN pin_475
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.00697211155331 100 82.25697211155331 ;
		END PORT
	END pin_475
	PIN pin_476
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.32669322709116 100 82.57669322709116 ;
		END PORT
	END pin_476
	PIN pin_477
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.646414342629 100 82.896414342629 ;
		END PORT
	END pin_477
	PIN pin_478
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.96613545816685 100 83.21613545816685 ;
		END PORT
	END pin_478
	PIN pin_479
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.28585657370469 100 83.53585657370469 ;
		END PORT
	END pin_479
	PIN pin_480
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.60557768924254 100 83.85557768924254 ;
		END PORT
	END pin_480
	PIN pin_481
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.92529880478038 100 84.17529880478038 ;
		END PORT
	END pin_481
	PIN pin_482
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.24501992031823 100 84.49501992031823 ;
		END PORT
	END pin_482
	PIN pin_483
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.56474103585607 100 84.81474103585607 ;
		END PORT
	END pin_483
	PIN pin_484
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.88446215139392 100 85.13446215139392 ;
		END PORT
	END pin_484
	PIN pin_485
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.20418326693176 100 85.45418326693176 ;
		END PORT
	END pin_485
	PIN pin_486
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.52390438246961 100 85.77390438246961 ;
		END PORT
	END pin_486
	PIN pin_487
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.84362549800746 100 86.09362549800746 ;
		END PORT
	END pin_487
	PIN pin_488
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.1633466135453 100 86.4133466135453 ;
		END PORT
	END pin_488
	PIN pin_489
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.48306772908315 100 86.73306772908315 ;
		END PORT
	END pin_489
	PIN pin_490
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.80278884462099 100 87.05278884462099 ;
		END PORT
	END pin_490
	PIN pin_491
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.12250996015884 100 87.37250996015884 ;
		END PORT
	END pin_491
	PIN pin_492
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.44223107569668 100 87.69223107569668 ;
		END PORT
	END pin_492
	PIN pin_493
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.76195219123453 100 88.01195219123453 ;
		END PORT
	END pin_493
	PIN pin_494
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.08167330677237 100 88.33167330677237 ;
		END PORT
	END pin_494
	PIN pin_495
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.40139442231022 100 88.65139442231022 ;
		END PORT
	END pin_495
	PIN pin_496
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.72111553784806 100 88.97111553784806 ;
		END PORT
	END pin_496
	PIN pin_497
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.04083665338591 100 89.29083665338591 ;
		END PORT
	END pin_497
	PIN pin_498
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.36055776892375 100 89.61055776892375 ;
		END PORT
	END pin_498
	PIN pin_499
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.6802788844616 100 89.9302788844616 ;
		END PORT
	END pin_499
	PIN pin_500
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.68027888446215 99.75 89.93027888446215 100 ;
		END PORT
	END pin_500
	PIN pin_501
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 89.36055776892431 99.75 89.61055776892431 100 ;
		END PORT
	END pin_501
	PIN pin_502
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.04083665338646 99.75 89.29083665338646 100 ;
		END PORT
	END pin_502
	PIN pin_503
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 88.72111553784862 99.75 88.97111553784862 100 ;
		END PORT
	END pin_503
	PIN pin_504
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.40139442231077 99.75 88.65139442231077 100 ;
		END PORT
	END pin_504
	PIN pin_505
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.08167330677293 99.75 88.33167330677293 100 ;
		END PORT
	END pin_505
	PIN pin_506
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.76195219123508 99.75 88.01195219123508 100 ;
		END PORT
	END pin_506
	PIN pin_507
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 87.44223107569724 99.75 87.69223107569724 100 ;
		END PORT
	END pin_507
	PIN pin_508
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.12250996015939 99.75 87.37250996015939 100 ;
		END PORT
	END pin_508
	PIN pin_509
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 86.80278884462155 99.75 87.05278884462155 100 ;
		END PORT
	END pin_509
	PIN pin_510
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.4830677290837 99.75 86.7330677290837 100 ;
		END PORT
	END pin_510
	PIN pin_511
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.16334661354585 99.75 86.41334661354585 100 ;
		END PORT
	END pin_511
	PIN pin_512
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 85.84362549800801 99.75 86.09362549800801 100 ;
		END PORT
	END pin_512
	PIN pin_513
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 85.52390438247016 99.75 85.77390438247016 100 ;
		END PORT
	END pin_513
	PIN pin_514
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.20418326693232 99.75 85.45418326693232 100 ;
		END PORT
	END pin_514
	PIN pin_515
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 84.88446215139447 99.75 85.13446215139447 100 ;
		END PORT
	END pin_515
	PIN pin_516
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 84.56474103585663 99.75 84.81474103585663 100 ;
		END PORT
	END pin_516
	PIN pin_517
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 84.24501992031878 99.75 84.49501992031878 100 ;
		END PORT
	END pin_517
	PIN pin_518
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 83.92529880478094 99.75 84.17529880478094 100 ;
		END PORT
	END pin_518
	PIN pin_519
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 83.60557768924309 99.75 83.85557768924309 100 ;
		END PORT
	END pin_519
	PIN pin_520
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.28585657370525 99.75 83.53585657370525 100 ;
		END PORT
	END pin_520
	PIN pin_521
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.9661354581674 99.75 83.2161354581674 100 ;
		END PORT
	END pin_521
	PIN pin_522
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.64641434262955 99.75 82.89641434262955 100 ;
		END PORT
	END pin_522
	PIN pin_523
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.32669322709171 99.75 82.57669322709171 100 ;
		END PORT
	END pin_523
	PIN pin_524
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.00697211155386 99.75 82.25697211155386 100 ;
		END PORT
	END pin_524
	PIN pin_525
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 81.68725099601602 99.75 81.93725099601602 100 ;
		END PORT
	END pin_525
	PIN pin_526
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.36752988047817 99.75 81.61752988047817 100 ;
		END PORT
	END pin_526
	PIN pin_527
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 81.04780876494033 99.75 81.29780876494033 100 ;
		END PORT
	END pin_527
	PIN pin_528
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 80.72808764940248 99.75 80.97808764940248 100 ;
		END PORT
	END pin_528
	PIN pin_529
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.40836653386464 99.75 80.65836653386464 100 ;
		END PORT
	END pin_529
	PIN pin_530
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 80.08864541832679 99.75 80.33864541832679 100 ;
		END PORT
	END pin_530
	PIN pin_531
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.76892430278895 99.75 80.01892430278895 100 ;
		END PORT
	END pin_531
	PIN pin_532
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 79.4492031872511 99.75 79.6992031872511 100 ;
		END PORT
	END pin_532
	PIN pin_533
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 79.12948207171326 99.75 79.37948207171326 100 ;
		END PORT
	END pin_533
	PIN pin_534
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 78.80976095617541 99.75 79.05976095617541 100 ;
		END PORT
	END pin_534
	PIN pin_535
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 78.49003984063756 99.75 78.74003984063756 100 ;
		END PORT
	END pin_535
	PIN pin_536
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 78.17031872509972 99.75 78.42031872509972 100 ;
		END PORT
	END pin_536
	PIN pin_537
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.85059760956187 99.75 78.10059760956187 100 ;
		END PORT
	END pin_537
	PIN pin_538
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.53087649402403 99.75 77.78087649402403 100 ;
		END PORT
	END pin_538
	PIN pin_539
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 77.21115537848618 99.75 77.46115537848618 100 ;
		END PORT
	END pin_539
	PIN pin_540
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 76.89143426294834 99.75 77.14143426294834 100 ;
		END PORT
	END pin_540
	PIN pin_541
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.57171314741049 99.75 76.82171314741049 100 ;
		END PORT
	END pin_541
	PIN pin_542
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.25199203187265 99.75 76.50199203187265 100 ;
		END PORT
	END pin_542
	PIN pin_543
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 75.9322709163348 99.75 76.1822709163348 100 ;
		END PORT
	END pin_543
	PIN pin_544
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 75.61254980079696 99.75 75.86254980079696 100 ;
		END PORT
	END pin_544
	PIN pin_545
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 75.29282868525911 99.75 75.54282868525911 100 ;
		END PORT
	END pin_545
	PIN pin_546
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 74.97310756972126 99.75 75.22310756972126 100 ;
		END PORT
	END pin_546
	PIN pin_547
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 74.65338645418342 99.75 74.90338645418342 100 ;
		END PORT
	END pin_547
	PIN pin_548
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 74.33366533864557 99.75 74.58366533864557 100 ;
		END PORT
	END pin_548
	PIN pin_549
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 74.01394422310773 99.75 74.26394422310773 100 ;
		END PORT
	END pin_549
	PIN pin_550
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 73.69422310756988 99.75 73.94422310756988 100 ;
		END PORT
	END pin_550
	PIN pin_551
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.37450199203204 99.75 73.62450199203204 100 ;
		END PORT
	END pin_551
	PIN pin_552
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.05478087649419 99.75 73.30478087649419 100 ;
		END PORT
	END pin_552
	PIN pin_553
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 72.73505976095635 99.75 72.98505976095635 100 ;
		END PORT
	END pin_553
	PIN pin_554
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 72.4153386454185 99.75 72.6653386454185 100 ;
		END PORT
	END pin_554
	PIN pin_555
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 72.09561752988066 99.75 72.34561752988066 100 ;
		END PORT
	END pin_555
	PIN pin_556
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 71.77589641434281 99.75 72.02589641434281 100 ;
		END PORT
	END pin_556
	PIN pin_557
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 71.45617529880496 99.75 71.70617529880496 100 ;
		END PORT
	END pin_557
	PIN pin_558
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 71.13645418326712 99.75 71.38645418326712 100 ;
		END PORT
	END pin_558
	PIN pin_559
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 70.81673306772927 99.75 71.06673306772927 100 ;
		END PORT
	END pin_559
	PIN pin_560
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.49701195219143 99.75 70.74701195219143 100 ;
		END PORT
	END pin_560
	PIN pin_561
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.17729083665358 99.75 70.42729083665358 100 ;
		END PORT
	END pin_561
	PIN pin_562
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 69.85756972111574 99.75 70.10756972111574 100 ;
		END PORT
	END pin_562
	PIN pin_563
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 69.53784860557789 99.75 69.78784860557789 100 ;
		END PORT
	END pin_563
	PIN pin_564
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 69.21812749004005 99.75 69.46812749004005 100 ;
		END PORT
	END pin_564
	PIN pin_565
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.8984063745022 99.75 69.1484063745022 100 ;
		END PORT
	END pin_565
	PIN pin_566
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 68.57868525896436 99.75 68.82868525896436 100 ;
		END PORT
	END pin_566
	PIN pin_567
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.25896414342651 99.75 68.50896414342651 100 ;
		END PORT
	END pin_567
	PIN pin_568
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 67.93924302788866 99.75 68.18924302788866 100 ;
		END PORT
	END pin_568
	PIN pin_569
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 67.61952191235082 99.75 67.86952191235082 100 ;
		END PORT
	END pin_569
	PIN pin_570
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.29980079681297 99.75 67.54980079681297 100 ;
		END PORT
	END pin_570
	PIN pin_571
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 66.98007968127513 99.75 67.23007968127513 100 ;
		END PORT
	END pin_571
	PIN pin_572
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.66035856573728 99.75 66.91035856573728 100 ;
		END PORT
	END pin_572
	PIN pin_573
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.34063745019944 99.75 66.59063745019944 100 ;
		END PORT
	END pin_573
	PIN pin_574
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.02091633466159 99.75 66.27091633466159 100 ;
		END PORT
	END pin_574
	PIN pin_575
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 65.70119521912375 99.75 65.95119521912375 100 ;
		END PORT
	END pin_575
	PIN pin_576
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 65.3814741035859 99.75 65.6314741035859 100 ;
		END PORT
	END pin_576
	PIN pin_577
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.06175298804806 99.75 65.31175298804806 100 ;
		END PORT
	END pin_577
	PIN pin_578
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.74203187251021 99.75 64.99203187251021 100 ;
		END PORT
	END pin_578
	PIN pin_579
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 64.42231075697237 99.75 64.67231075697237 100 ;
		END PORT
	END pin_579
	PIN pin_580
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 64.10258964143452 99.75 64.35258964143452 100 ;
		END PORT
	END pin_580
	PIN pin_581
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.782868525896674 99.75 64.03286852589667 100 ;
		END PORT
	END pin_581
	PIN pin_582
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.46314741035883 99.75 63.71314741035883 100 ;
		END PORT
	END pin_582
	PIN pin_583
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 63.14342629482098 99.75 63.39342629482098 100 ;
		END PORT
	END pin_583
	PIN pin_584
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.82370517928314 99.75 63.07370517928314 100 ;
		END PORT
	END pin_584
	PIN pin_585
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.50398406374529 99.75 62.75398406374529 100 ;
		END PORT
	END pin_585
	PIN pin_586
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 62.18426294820745 99.75 62.43426294820745 100 ;
		END PORT
	END pin_586
	PIN pin_587
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 61.8645418326696 99.75 62.1145418326696 100 ;
		END PORT
	END pin_587
	PIN pin_588
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 61.544820717131756 99.75 61.794820717131756 100 ;
		END PORT
	END pin_588
	PIN pin_589
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 61.22509960159391 99.75 61.47509960159391 100 ;
		END PORT
	END pin_589
	PIN pin_590
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 60.905378486056065 99.75 61.155378486056065 100 ;
		END PORT
	END pin_590
	PIN pin_591
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 60.58565737051822 99.75 60.83565737051822 100 ;
		END PORT
	END pin_591
	PIN pin_592
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 60.265936254980375 99.75 60.515936254980375 100 ;
		END PORT
	END pin_592
	PIN pin_593
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 59.94621513944253 99.75 60.19621513944253 100 ;
		END PORT
	END pin_593
	PIN pin_594
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 59.626494023904684 99.75 59.876494023904684 100 ;
		END PORT
	END pin_594
	PIN pin_595
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 59.30677290836684 99.75 59.55677290836684 100 ;
		END PORT
	END pin_595
	PIN pin_596
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.98705179282899 99.75 59.23705179282899 100 ;
		END PORT
	END pin_596
	PIN pin_597
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.66733067729115 99.75 58.91733067729115 100 ;
		END PORT
	END pin_597
	PIN pin_598
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.3476095617533 99.75 58.5976095617533 100 ;
		END PORT
	END pin_598
	PIN pin_599
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.02788844621546 99.75 58.27788844621546 100 ;
		END PORT
	END pin_599
	PIN pin_600
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.70816733067761 99.75 57.95816733067761 100 ;
		END PORT
	END pin_600
	PIN pin_601
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 57.388446215139766 99.75 57.638446215139766 100 ;
		END PORT
	END pin_601
	PIN pin_602
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 57.06872509960192 99.75 57.31872509960192 100 ;
		END PORT
	END pin_602
	PIN pin_603
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.749003984064075 99.75 56.999003984064075 100 ;
		END PORT
	END pin_603
	PIN pin_604
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.42928286852623 99.75 56.67928286852623 100 ;
		END PORT
	END pin_604
	PIN pin_605
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.109561752988384 99.75 56.359561752988384 100 ;
		END PORT
	END pin_605
	PIN pin_606
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 55.78984063745054 99.75 56.03984063745054 100 ;
		END PORT
	END pin_606
	PIN pin_607
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 55.47011952191269 99.75 55.72011952191269 100 ;
		END PORT
	END pin_607
	PIN pin_608
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.15039840637485 99.75 55.40039840637485 100 ;
		END PORT
	END pin_608
	PIN pin_609
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 54.830677290837 99.75 55.080677290837 100 ;
		END PORT
	END pin_609
	PIN pin_610
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 54.51095617529916 99.75 54.76095617529916 100 ;
		END PORT
	END pin_610
	PIN pin_611
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 54.19123505976131 99.75 54.44123505976131 100 ;
		END PORT
	END pin_611
	PIN pin_612
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 53.871513944223466 99.75 54.121513944223466 100 ;
		END PORT
	END pin_612
	PIN pin_613
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 53.55179282868562 99.75 53.80179282868562 100 ;
		END PORT
	END pin_613
	PIN pin_614
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.232071713147775 99.75 53.482071713147775 100 ;
		END PORT
	END pin_614
	PIN pin_615
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 52.91235059760993 99.75 53.16235059760993 100 ;
		END PORT
	END pin_615
	PIN pin_616
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 52.592629482072084 99.75 52.842629482072084 100 ;
		END PORT
	END pin_616
	PIN pin_617
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 52.27290836653424 99.75 52.52290836653424 100 ;
		END PORT
	END pin_617
	PIN pin_618
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 51.95318725099639 99.75 52.20318725099639 100 ;
		END PORT
	END pin_618
	PIN pin_619
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.63346613545855 99.75 51.88346613545855 100 ;
		END PORT
	END pin_619
	PIN pin_620
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 51.3137450199207 99.75 51.5637450199207 100 ;
		END PORT
	END pin_620
	PIN pin_621
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 50.99402390438286 99.75 51.24402390438286 100 ;
		END PORT
	END pin_621
	PIN pin_622
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.67430278884501 99.75 50.92430278884501 100 ;
		END PORT
	END pin_622
	PIN pin_623
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.354581673307166 99.75 50.604581673307166 100 ;
		END PORT
	END pin_623
	PIN pin_624
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.03486055776932 99.75 50.28486055776932 100 ;
		END PORT
	END pin_624
	PIN pin_625
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 49.715139442231475 99.75 49.965139442231475 100 ;
		END PORT
	END pin_625
	PIN pin_626
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 49.39541832669363 99.75 49.64541832669363 100 ;
		END PORT
	END pin_626
	PIN pin_627
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 49.075697211155784 99.75 49.325697211155784 100 ;
		END PORT
	END pin_627
	PIN pin_628
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 48.75597609561794 99.75 49.00597609561794 100 ;
		END PORT
	END pin_628
	PIN pin_629
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 48.43625498008009 99.75 48.68625498008009 100 ;
		END PORT
	END pin_629
	PIN pin_630
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.11653386454225 99.75 48.36653386454225 100 ;
		END PORT
	END pin_630
	PIN pin_631
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.7968127490044 99.75 48.0468127490044 100 ;
		END PORT
	END pin_631
	PIN pin_632
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 47.47709163346656 99.75 47.72709163346656 100 ;
		END PORT
	END pin_632
	PIN pin_633
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.15737051792871 99.75 47.40737051792871 100 ;
		END PORT
	END pin_633
	PIN pin_634
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 46.837649402390866 99.75 47.087649402390866 100 ;
		END PORT
	END pin_634
	PIN pin_635
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 46.51792828685302 99.75 46.76792828685302 100 ;
		END PORT
	END pin_635
	PIN pin_636
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.198207171315175 99.75 46.448207171315175 100 ;
		END PORT
	END pin_636
	PIN pin_637
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 45.87848605577733 99.75 46.12848605577733 100 ;
		END PORT
	END pin_637
	PIN pin_638
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.558764940239485 99.75 45.808764940239485 100 ;
		END PORT
	END pin_638
	PIN pin_639
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.23904382470164 99.75 45.48904382470164 100 ;
		END PORT
	END pin_639
	PIN pin_640
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 44.919322709163794 99.75 45.169322709163794 100 ;
		END PORT
	END pin_640
	PIN pin_641
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.59960159362595 99.75 44.84960159362595 100 ;
		END PORT
	END pin_641
	PIN pin_642
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 44.2798804780881 99.75 44.5298804780881 100 ;
		END PORT
	END pin_642
	PIN pin_643
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.96015936255026 99.75 44.21015936255026 100 ;
		END PORT
	END pin_643
	PIN pin_644
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.64043824701241 99.75 43.89043824701241 100 ;
		END PORT
	END pin_644
	PIN pin_645
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.32071713147457 99.75 43.57071713147457 100 ;
		END PORT
	END pin_645
	PIN pin_646
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.00099601593672 99.75 43.25099601593672 100 ;
		END PORT
	END pin_646
	PIN pin_647
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 42.681274900398876 99.75 42.931274900398876 100 ;
		END PORT
	END pin_647
	PIN pin_648
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.36155378486103 99.75 42.61155378486103 100 ;
		END PORT
	END pin_648
	PIN pin_649
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 42.041832669323185 99.75 42.291832669323185 100 ;
		END PORT
	END pin_649
	PIN pin_650
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 41.72211155378534 99.75 41.97211155378534 100 ;
		END PORT
	END pin_650
	PIN pin_651
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 41.402390438247494 99.75 41.652390438247494 100 ;
		END PORT
	END pin_651
	PIN pin_652
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.08266932270965 99.75 41.33266932270965 100 ;
		END PORT
	END pin_652
	PIN pin_653
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 40.7629482071718 99.75 41.0129482071718 100 ;
		END PORT
	END pin_653
	PIN pin_654
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.44322709163396 99.75 40.69322709163396 100 ;
		END PORT
	END pin_654
	PIN pin_655
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 40.12350597609611 99.75 40.37350597609611 100 ;
		END PORT
	END pin_655
	PIN pin_656
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 39.80378486055827 99.75 40.05378486055827 100 ;
		END PORT
	END pin_656
	PIN pin_657
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 39.48406374502042 99.75 39.73406374502042 100 ;
		END PORT
	END pin_657
	PIN pin_658
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 39.164342629482576 99.75 39.414342629482576 100 ;
		END PORT
	END pin_658
	PIN pin_659
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.84462151394473 99.75 39.09462151394473 100 ;
		END PORT
	END pin_659
	PIN pin_660
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 38.524900398406885 99.75 38.774900398406885 100 ;
		END PORT
	END pin_660
	PIN pin_661
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.20517928286904 99.75 38.45517928286904 100 ;
		END PORT
	END pin_661
	PIN pin_662
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 37.885458167331194 99.75 38.135458167331194 100 ;
		END PORT
	END pin_662
	PIN pin_663
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.56573705179335 99.75 37.81573705179335 100 ;
		END PORT
	END pin_663
	PIN pin_664
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 37.2460159362555 99.75 37.4960159362555 100 ;
		END PORT
	END pin_664
	PIN pin_665
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 36.92629482071766 99.75 37.17629482071766 100 ;
		END PORT
	END pin_665
	PIN pin_666
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 36.60657370517981 99.75 36.85657370517981 100 ;
		END PORT
	END pin_666
	PIN pin_667
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.28685258964197 99.75 36.53685258964197 100 ;
		END PORT
	END pin_667
	PIN pin_668
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 35.96713147410412 99.75 36.21713147410412 100 ;
		END PORT
	END pin_668
	PIN pin_669
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 35.647410358566276 99.75 35.897410358566276 100 ;
		END PORT
	END pin_669
	PIN pin_670
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.32768924302843 99.75 35.57768924302843 100 ;
		END PORT
	END pin_670
	PIN pin_671
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.007968127490585 99.75 35.257968127490585 100 ;
		END PORT
	END pin_671
	PIN pin_672
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 34.68824701195274 99.75 34.93824701195274 100 ;
		END PORT
	END pin_672
	PIN pin_673
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.368525896414894 99.75 34.618525896414894 100 ;
		END PORT
	END pin_673
	PIN pin_674
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 34.04880478087705 99.75 34.29880478087705 100 ;
		END PORT
	END pin_674
	PIN pin_675
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.7290836653392 99.75 33.9790836653392 100 ;
		END PORT
	END pin_675
	PIN pin_676
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 33.40936254980136 99.75 33.65936254980136 100 ;
		END PORT
	END pin_676
	PIN pin_677
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.08964143426351 99.75 33.33964143426351 100 ;
		END PORT
	END pin_677
	PIN pin_678
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.76992031872567 99.75 33.01992031872567 100 ;
		END PORT
	END pin_678
	PIN pin_679
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.45019920318782 99.75 32.70019920318782 100 ;
		END PORT
	END pin_679
	PIN pin_680
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 32.130478087649976 99.75 32.380478087649976 100 ;
		END PORT
	END pin_680
	PIN pin_681
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.81075697211213 99.75 32.06075697211213 100 ;
		END PORT
	END pin_681
	PIN pin_682
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 31.491035856574282 99.75 31.741035856574282 100 ;
		END PORT
	END pin_682
	PIN pin_683
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.171314741036433 99.75 31.421314741036433 100 ;
		END PORT
	END pin_683
	PIN pin_684
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 30.851593625498584 99.75 31.101593625498584 100 ;
		END PORT
	END pin_684
	PIN pin_685
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 30.531872509960735 99.75 30.781872509960735 100 ;
		END PORT
	END pin_685
	PIN pin_686
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 30.212151394422886 99.75 30.462151394422886 100 ;
		END PORT
	END pin_686
	PIN pin_687
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.892430278885037 99.75 30.142430278885037 100 ;
		END PORT
	END pin_687
	PIN pin_688
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.572709163347188 99.75 29.822709163347188 100 ;
		END PORT
	END pin_688
	PIN pin_689
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.25298804780934 99.75 29.50298804780934 100 ;
		END PORT
	END pin_689
	PIN pin_690
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.93326693227149 99.75 29.18326693227149 100 ;
		END PORT
	END pin_690
	PIN pin_691
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 28.61354581673364 99.75 28.86354581673364 100 ;
		END PORT
	END pin_691
	PIN pin_692
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 28.293824701195792 99.75 28.543824701195792 100 ;
		END PORT
	END pin_692
	PIN pin_693
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.974103585657943 99.75 28.224103585657943 100 ;
		END PORT
	END pin_693
	PIN pin_694
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.654382470120094 99.75 27.904382470120094 100 ;
		END PORT
	END pin_694
	PIN pin_695
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 27.334661354582245 99.75 27.584661354582245 100 ;
		END PORT
	END pin_695
	PIN pin_696
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.014940239044396 99.75 27.264940239044396 100 ;
		END PORT
	END pin_696
	PIN pin_697
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 26.695219123506547 99.75 26.945219123506547 100 ;
		END PORT
	END pin_697
	PIN pin_698
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.375498007968698 99.75 26.625498007968698 100 ;
		END PORT
	END pin_698
	PIN pin_699
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.05577689243085 99.75 26.30577689243085 100 ;
		END PORT
	END pin_699
	PIN pin_700
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 25.736055776893 99.75 25.986055776893 100 ;
		END PORT
	END pin_700
	PIN pin_701
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 25.41633466135515 99.75 25.66633466135515 100 ;
		END PORT
	END pin_701
	PIN pin_702
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 25.096613545817302 99.75 25.346613545817302 100 ;
		END PORT
	END pin_702
	PIN pin_703
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.776892430279453 99.75 25.026892430279453 100 ;
		END PORT
	END pin_703
	PIN pin_704
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 24.457171314741604 99.75 24.707171314741604 100 ;
		END PORT
	END pin_704
	PIN pin_705
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.137450199203755 99.75 24.387450199203755 100 ;
		END PORT
	END pin_705
	PIN pin_706
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.817729083665906 99.75 24.067729083665906 100 ;
		END PORT
	END pin_706
	PIN pin_707
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 23.498007968128057 99.75 23.748007968128057 100 ;
		END PORT
	END pin_707
	PIN pin_708
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 23.178286852590208 99.75 23.428286852590208 100 ;
		END PORT
	END pin_708
	PIN pin_709
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.85856573705236 99.75 23.10856573705236 100 ;
		END PORT
	END pin_709
	PIN pin_710
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 22.53884462151451 99.75 22.78884462151451 100 ;
		END PORT
	END pin_710
	PIN pin_711
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.21912350597666 99.75 22.46912350597666 100 ;
		END PORT
	END pin_711
	PIN pin_712
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 21.899402390438812 99.75 22.149402390438812 100 ;
		END PORT
	END pin_712
	PIN pin_713
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 21.579681274900963 99.75 21.829681274900963 100 ;
		END PORT
	END pin_713
	PIN pin_714
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 21.259960159363114 99.75 21.509960159363114 100 ;
		END PORT
	END pin_714
	PIN pin_715
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.940239043825265 99.75 21.190239043825265 100 ;
		END PORT
	END pin_715
	PIN pin_716
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.620517928287416 99.75 20.870517928287416 100 ;
		END PORT
	END pin_716
	PIN pin_717
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 20.300796812749567 99.75 20.550796812749567 100 ;
		END PORT
	END pin_717
	PIN pin_718
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 19.98107569721172 99.75 20.23107569721172 100 ;
		END PORT
	END pin_718
	PIN pin_719
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.66135458167387 99.75 19.91135458167387 100 ;
		END PORT
	END pin_719
	PIN pin_720
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.34163346613602 99.75 19.59163346613602 100 ;
		END PORT
	END pin_720
	PIN pin_721
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.02191235059817 99.75 19.27191235059817 100 ;
		END PORT
	END pin_721
	PIN pin_722
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 18.702191235060322 99.75 18.952191235060322 100 ;
		END PORT
	END pin_722
	PIN pin_723
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.382470119522473 99.75 18.632470119522473 100 ;
		END PORT
	END pin_723
	PIN pin_724
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 18.062749003984624 99.75 18.312749003984624 100 ;
		END PORT
	END pin_724
	PIN pin_725
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 17.743027888446775 99.75 17.993027888446775 100 ;
		END PORT
	END pin_725
	PIN pin_726
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 17.423306772908926 99.75 17.673306772908926 100 ;
		END PORT
	END pin_726
	PIN pin_727
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.103585657371077 99.75 17.353585657371077 100 ;
		END PORT
	END pin_727
	PIN pin_728
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 16.78386454183323 99.75 17.03386454183323 100 ;
		END PORT
	END pin_728
	PIN pin_729
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.46414342629538 99.75 16.71414342629538 100 ;
		END PORT
	END pin_729
	PIN pin_730
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.14442231075753 99.75 16.39442231075753 100 ;
		END PORT
	END pin_730
	PIN pin_731
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.824701195219681 99.75 16.07470119521968 100 ;
		END PORT
	END pin_731
	PIN pin_732
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.504980079681832 99.75 15.754980079681832 100 ;
		END PORT
	END pin_732
	PIN pin_733
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.185258964143983 99.75 15.435258964143983 100 ;
		END PORT
	END pin_733
	PIN pin_734
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 14.865537848606134 99.75 15.115537848606134 100 ;
		END PORT
	END pin_734
	PIN pin_735
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 14.545816733068285 99.75 14.795816733068285 100 ;
		END PORT
	END pin_735
	PIN pin_736
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 14.226095617530436 99.75 14.476095617530436 100 ;
		END PORT
	END pin_736
	PIN pin_737
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 13.906374501992588 99.75 14.156374501992588 100 ;
		END PORT
	END pin_737
	PIN pin_738
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 13.586653386454739 99.75 13.836653386454739 100 ;
		END PORT
	END pin_738
	PIN pin_739
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 13.26693227091689 99.75 13.51693227091689 100 ;
		END PORT
	END pin_739
	PIN pin_740
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 12.94721115537904 99.75 13.19721115537904 100 ;
		END PORT
	END pin_740
	PIN pin_741
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 12.627490039841192 99.75 12.877490039841192 100 ;
		END PORT
	END pin_741
	PIN pin_742
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 12.307768924303343 99.75 12.557768924303343 100 ;
		END PORT
	END pin_742
	PIN pin_743
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.988047808765494 99.75 12.238047808765494 100 ;
		END PORT
	END pin_743
	PIN pin_744
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.668326693227645 99.75 11.918326693227645 100 ;
		END PORT
	END pin_744
	PIN pin_745
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 11.348605577689796 99.75 11.598605577689796 100 ;
		END PORT
	END pin_745
	PIN pin_746
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.028884462151947 99.75 11.278884462151947 100 ;
		END PORT
	END pin_746
	PIN pin_747
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 10.709163346614098 99.75 10.959163346614098 100 ;
		END PORT
	END pin_747
	PIN pin_748
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 10.389442231076249 99.75 10.639442231076249 100 ;
		END PORT
	END pin_748
	PIN pin_749
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 10.0697211155384 99.75 10.3197211155384 100 ;
		END PORT
	END pin_749
	PIN pin_750
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 10.069721115537849 0 10.319721115537849 0.25 ;
		END PORT
	END pin_750
	PIN pin_751
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 10.389442231075698 0 10.639442231075698 0.25 ;
		END PORT
	END pin_751
	PIN pin_752
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 10.709163346613547 0 10.959163346613547 0.25 ;
		END PORT
	END pin_752
	PIN pin_753
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 11.028884462151396 0 11.278884462151396 0.25 ;
		END PORT
	END pin_753
	PIN pin_754
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.348605577689245 0 11.598605577689245 0.25 ;
		END PORT
	END pin_754
	PIN pin_755
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.668326693227094 0 11.918326693227094 0.25 ;
		END PORT
	END pin_755
	PIN pin_756
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.988047808764943 0 12.238047808764943 0.25 ;
		END PORT
	END pin_756
	PIN pin_757
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 12.307768924302792 0 12.557768924302792 0.25 ;
		END PORT
	END pin_757
	PIN pin_758
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 12.627490039840641 0 12.877490039840641 0.25 ;
		END PORT
	END pin_758
	PIN pin_759
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 12.94721115537849 0 13.19721115537849 0.25 ;
		END PORT
	END pin_759
	PIN pin_760
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 13.266932270916339 0 13.516932270916339 0.25 ;
		END PORT
	END pin_760
	PIN pin_761
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 13.586653386454188 0 13.836653386454188 0.25 ;
		END PORT
	END pin_761
	PIN pin_762
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 13.906374501992037 0 14.156374501992037 0.25 ;
		END PORT
	END pin_762
	PIN pin_763
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 14.226095617529886 0 14.476095617529886 0.25 ;
		END PORT
	END pin_763
	PIN pin_764
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.545816733067735 0 14.795816733067735 0.25 ;
		END PORT
	END pin_764
	PIN pin_765
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.865537848605584 0 15.115537848605584 0.25 ;
		END PORT
	END pin_765
	PIN pin_766
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.185258964143433 0 15.435258964143433 0.25 ;
		END PORT
	END pin_766
	PIN pin_767
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.504980079681282 0 15.754980079681282 0.25 ;
		END PORT
	END pin_767
	PIN pin_768
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.82470119521913 0 16.07470119521913 0.25 ;
		END PORT
	END pin_768
	PIN pin_769
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.14442231075698 0 16.39442231075698 0.25 ;
		END PORT
	END pin_769
	PIN pin_770
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 16.46414342629483 0 16.71414342629483 0.25 ;
		END PORT
	END pin_770
	PIN pin_771
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.783864541832678 0 17.033864541832678 0.25 ;
		END PORT
	END pin_771
	PIN pin_772
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 17.103585657370527 0 17.353585657370527 0.25 ;
		END PORT
	END pin_772
	PIN pin_773
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 17.423306772908376 0 17.673306772908376 0.25 ;
		END PORT
	END pin_773
	PIN pin_774
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 17.743027888446225 0 17.993027888446225 0.25 ;
		END PORT
	END pin_774
	PIN pin_775
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 18.062749003984074 0 18.312749003984074 0.25 ;
		END PORT
	END pin_775
	PIN pin_776
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.382470119521923 0 18.632470119521923 0.25 ;
		END PORT
	END pin_776
	PIN pin_777
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.70219123505977 0 18.95219123505977 0.25 ;
		END PORT
	END pin_777
	PIN pin_778
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.02191235059762 0 19.27191235059762 0.25 ;
		END PORT
	END pin_778
	PIN pin_779
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.34163346613547 0 19.59163346613547 0.25 ;
		END PORT
	END pin_779
	PIN pin_780
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.66135458167332 0 19.91135458167332 0.25 ;
		END PORT
	END pin_780
	PIN pin_781
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 19.981075697211168 0 20.231075697211168 0.25 ;
		END PORT
	END pin_781
	PIN pin_782
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.300796812749017 0 20.550796812749017 0.25 ;
		END PORT
	END pin_782
	PIN pin_783
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 20.620517928286866 0 20.870517928286866 0.25 ;
		END PORT
	END pin_783
	PIN pin_784
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 20.940239043824715 0 21.190239043824715 0.25 ;
		END PORT
	END pin_784
	PIN pin_785
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.259960159362564 0 21.509960159362564 0.25 ;
		END PORT
	END pin_785
	PIN pin_786
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.579681274900413 0 21.829681274900413 0.25 ;
		END PORT
	END pin_786
	PIN pin_787
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 21.89940239043826 0 22.14940239043826 0.25 ;
		END PORT
	END pin_787
	PIN pin_788
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.21912350597611 0 22.46912350597611 0.25 ;
		END PORT
	END pin_788
	PIN pin_789
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.53884462151396 0 22.78884462151396 0.25 ;
		END PORT
	END pin_789
	PIN pin_790
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.85856573705181 0 23.10856573705181 0.25 ;
		END PORT
	END pin_790
	PIN pin_791
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.178286852589657 0 23.428286852589657 0.25 ;
		END PORT
	END pin_791
	PIN pin_792
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 23.498007968127506 0 23.748007968127506 0.25 ;
		END PORT
	END pin_792
	PIN pin_793
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.817729083665355 0 24.067729083665355 0.25 ;
		END PORT
	END pin_793
	PIN pin_794
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 24.137450199203204 0 24.387450199203204 0.25 ;
		END PORT
	END pin_794
	PIN pin_795
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.457171314741053 0 24.707171314741053 0.25 ;
		END PORT
	END pin_795
	PIN pin_796
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.776892430278902 0 25.026892430278902 0.25 ;
		END PORT
	END pin_796
	PIN pin_797
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 25.09661354581675 0 25.34661354581675 0.25 ;
		END PORT
	END pin_797
	PIN pin_798
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 25.4163346613546 0 25.6663346613546 0.25 ;
		END PORT
	END pin_798
	PIN pin_799
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 25.73605577689245 0 25.98605577689245 0.25 ;
		END PORT
	END pin_799
	PIN pin_800
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 26.0557768924303 0 26.3057768924303 0.25 ;
		END PORT
	END pin_800
	PIN pin_801
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.375498007968147 0 26.625498007968147 0.25 ;
		END PORT
	END pin_801
	PIN pin_802
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.695219123505996 0 26.945219123505996 0.25 ;
		END PORT
	END pin_802
	PIN pin_803
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.014940239043845 0 27.264940239043845 0.25 ;
		END PORT
	END pin_803
	PIN pin_804
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.334661354581694 0 27.584661354581694 0.25 ;
		END PORT
	END pin_804
	PIN pin_805
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.654382470119543 0 27.904382470119543 0.25 ;
		END PORT
	END pin_805
	PIN pin_806
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 27.974103585657392 0 28.224103585657392 0.25 ;
		END PORT
	END pin_806
	PIN pin_807
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 28.29382470119524 0 28.54382470119524 0.25 ;
		END PORT
	END pin_807
	PIN pin_808
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.61354581673309 0 28.86354581673309 0.25 ;
		END PORT
	END pin_808
	PIN pin_809
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 28.93326693227094 0 29.18326693227094 0.25 ;
		END PORT
	END pin_809
	PIN pin_810
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.25298804780879 0 29.50298804780879 0.25 ;
		END PORT
	END pin_810
	PIN pin_811
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 29.572709163346637 0 29.822709163346637 0.25 ;
		END PORT
	END pin_811
	PIN pin_812
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.892430278884486 0 30.142430278884486 0.25 ;
		END PORT
	END pin_812
	PIN pin_813
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.212151394422335 0 30.462151394422335 0.25 ;
		END PORT
	END pin_813
	PIN pin_814
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 30.531872509960184 0 30.781872509960184 0.25 ;
		END PORT
	END pin_814
	PIN pin_815
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.851593625498033 0 31.101593625498033 0.25 ;
		END PORT
	END pin_815
	PIN pin_816
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 31.171314741035882 0 31.421314741035882 0.25 ;
		END PORT
	END pin_816
	PIN pin_817
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.49103585657373 0 31.74103585657373 0.25 ;
		END PORT
	END pin_817
	PIN pin_818
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.81075697211158 0 32.06075697211158 0.25 ;
		END PORT
	END pin_818
	PIN pin_819
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.13047808764942 0 32.38047808764942 0.25 ;
		END PORT
	END pin_819
	PIN pin_820
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 32.45019920318727 0 32.70019920318727 0.25 ;
		END PORT
	END pin_820
	PIN pin_821
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 32.76992031872511 0 33.01992031872511 0.25 ;
		END PORT
	END pin_821
	PIN pin_822
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 33.08964143426296 0 33.33964143426296 0.25 ;
		END PORT
	END pin_822
	PIN pin_823
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.409362549800804 0 33.659362549800804 0.25 ;
		END PORT
	END pin_823
	PIN pin_824
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 33.72908366533865 0 33.97908366533865 0.25 ;
		END PORT
	END pin_824
	PIN pin_825
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 34.048804780876495 0 34.298804780876495 0.25 ;
		END PORT
	END pin_825
	PIN pin_826
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.36852589641434 0 34.61852589641434 0.25 ;
		END PORT
	END pin_826
	PIN pin_827
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 34.688247011952186 0 34.938247011952186 0.25 ;
		END PORT
	END pin_827
	PIN pin_828
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.00796812749003 0 35.25796812749003 0.25 ;
		END PORT
	END pin_828
	PIN pin_829
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 35.327689243027876 0 35.577689243027876 0.25 ;
		END PORT
	END pin_829
	PIN pin_830
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.64741035856572 0 35.89741035856572 0.25 ;
		END PORT
	END pin_830
	PIN pin_831
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.96713147410357 0 36.21713147410357 0.25 ;
		END PORT
	END pin_831
	PIN pin_832
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 36.28685258964141 0 36.53685258964141 0.25 ;
		END PORT
	END pin_832
	PIN pin_833
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.60657370517926 0 36.85657370517926 0.25 ;
		END PORT
	END pin_833
	PIN pin_834
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.926294820717104 0 37.176294820717104 0.25 ;
		END PORT
	END pin_834
	PIN pin_835
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.24601593625495 0 37.49601593625495 0.25 ;
		END PORT
	END pin_835
	PIN pin_836
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 37.565737051792794 0 37.815737051792794 0.25 ;
		END PORT
	END pin_836
	PIN pin_837
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.88545816733064 0 38.13545816733064 0.25 ;
		END PORT
	END pin_837
	PIN pin_838
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.205179282868485 0 38.455179282868485 0.25 ;
		END PORT
	END pin_838
	PIN pin_839
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.52490039840633 0 38.77490039840633 0.25 ;
		END PORT
	END pin_839
	PIN pin_840
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 38.844621513944176 0 39.094621513944176 0.25 ;
		END PORT
	END pin_840
	PIN pin_841
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 39.16434262948202 0 39.41434262948202 0.25 ;
		END PORT
	END pin_841
	PIN pin_842
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 39.48406374501987 0 39.73406374501987 0.25 ;
		END PORT
	END pin_842
	PIN pin_843
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 39.80378486055771 0 40.05378486055771 0.25 ;
		END PORT
	END pin_843
	PIN pin_844
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 40.12350597609556 0 40.37350597609556 0.25 ;
		END PORT
	END pin_844
	PIN pin_845
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 40.4432270916334 0 40.6932270916334 0.25 ;
		END PORT
	END pin_845
	PIN pin_846
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 40.76294820717125 0 41.01294820717125 0.25 ;
		END PORT
	END pin_846
	PIN pin_847
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.082669322709094 0 41.332669322709094 0.25 ;
		END PORT
	END pin_847
	PIN pin_848
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.40239043824694 0 41.65239043824694 0.25 ;
		END PORT
	END pin_848
	PIN pin_849
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 41.722111553784785 0 41.972111553784785 0.25 ;
		END PORT
	END pin_849
	PIN pin_850
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.04183266932263 0 42.29183266932263 0.25 ;
		END PORT
	END pin_850
	PIN pin_851
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 42.361553784860476 0 42.611553784860476 0.25 ;
		END PORT
	END pin_851
	PIN pin_852
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.68127490039832 0 42.93127490039832 0.25 ;
		END PORT
	END pin_852
	PIN pin_853
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.00099601593617 0 43.25099601593617 0.25 ;
		END PORT
	END pin_853
	PIN pin_854
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 43.32071713147401 0 43.57071713147401 0.25 ;
		END PORT
	END pin_854
	PIN pin_855
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.64043824701186 0 43.89043824701186 0.25 ;
		END PORT
	END pin_855
	PIN pin_856
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.9601593625497 0 44.2101593625497 0.25 ;
		END PORT
	END pin_856
	PIN pin_857
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 44.27988047808755 0 44.52988047808755 0.25 ;
		END PORT
	END pin_857
	PIN pin_858
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 44.599601593625394 0 44.849601593625394 0.25 ;
		END PORT
	END pin_858
	PIN pin_859
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.91932270916324 0 45.16932270916324 0.25 ;
		END PORT
	END pin_859
	PIN pin_860
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 45.239043824701085 0 45.489043824701085 0.25 ;
		END PORT
	END pin_860
	PIN pin_861
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.55876494023893 0 45.80876494023893 0.25 ;
		END PORT
	END pin_861
	PIN pin_862
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 45.878486055776776 0 46.128486055776776 0.25 ;
		END PORT
	END pin_862
	PIN pin_863
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.19820717131462 0 46.44820717131462 0.25 ;
		END PORT
	END pin_863
	PIN pin_864
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.51792828685247 0 46.76792828685247 0.25 ;
		END PORT
	END pin_864
	PIN pin_865
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 46.83764940239031 0 47.08764940239031 0.25 ;
		END PORT
	END pin_865
	PIN pin_866
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.15737051792816 0 47.40737051792816 0.25 ;
		END PORT
	END pin_866
	PIN pin_867
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 47.477091633466 0 47.727091633466 0.25 ;
		END PORT
	END pin_867
	PIN pin_868
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.79681274900385 0 48.04681274900385 0.25 ;
		END PORT
	END pin_868
	PIN pin_869
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 48.116533864541694 0 48.366533864541694 0.25 ;
		END PORT
	END pin_869
	PIN pin_870
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.43625498007954 0 48.68625498007954 0.25 ;
		END PORT
	END pin_870
	PIN pin_871
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 48.755976095617385 0 49.005976095617385 0.25 ;
		END PORT
	END pin_871
	PIN pin_872
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.07569721115523 0 49.32569721115523 0.25 ;
		END PORT
	END pin_872
	PIN pin_873
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 49.395418326693076 0 49.645418326693076 0.25 ;
		END PORT
	END pin_873
	PIN pin_874
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 49.71513944223092 0 49.96513944223092 0.25 ;
		END PORT
	END pin_874
	PIN pin_875
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.034860557768766 0 50.284860557768766 0.25 ;
		END PORT
	END pin_875
	PIN pin_876
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.35458167330661 0 50.60458167330661 0.25 ;
		END PORT
	END pin_876
	PIN pin_877
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 50.67430278884446 0 50.92430278884446 0.25 ;
		END PORT
	END pin_877
	PIN pin_878
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 50.9940239043823 0 51.2440239043823 0.25 ;
		END PORT
	END pin_878
	PIN pin_879
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.31374501992015 0 51.56374501992015 0.25 ;
		END PORT
	END pin_879
	PIN pin_880
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 51.633466135457994 0 51.883466135457994 0.25 ;
		END PORT
	END pin_880
	PIN pin_881
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.95318725099584 0 52.20318725099584 0.25 ;
		END PORT
	END pin_881
	PIN pin_882
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 52.272908366533684 0 52.522908366533684 0.25 ;
		END PORT
	END pin_882
	PIN pin_883
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 52.59262948207153 0 52.84262948207153 0.25 ;
		END PORT
	END pin_883
	PIN pin_884
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 52.912350597609375 0 53.162350597609375 0.25 ;
		END PORT
	END pin_884
	PIN pin_885
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 53.23207171314722 0 53.48207171314722 0.25 ;
		END PORT
	END pin_885
	PIN pin_886
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.551792828685066 0 53.801792828685066 0.25 ;
		END PORT
	END pin_886
	PIN pin_887
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.87151394422291 0 54.12151394422291 0.25 ;
		END PORT
	END pin_887
	PIN pin_888
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 54.19123505976076 0 54.44123505976076 0.25 ;
		END PORT
	END pin_888
	PIN pin_889
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 54.5109561752986 0 54.7609561752986 0.25 ;
		END PORT
	END pin_889
	PIN pin_890
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 54.83067729083645 0 55.08067729083645 0.25 ;
		END PORT
	END pin_890
	PIN pin_891
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 55.15039840637429 0 55.40039840637429 0.25 ;
		END PORT
	END pin_891
	PIN pin_892
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 55.47011952191214 0 55.72011952191214 0.25 ;
		END PORT
	END pin_892
	PIN pin_893
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.789840637449984 0 56.039840637449984 0.25 ;
		END PORT
	END pin_893
	PIN pin_894
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.10956175298783 0 56.35956175298783 0.25 ;
		END PORT
	END pin_894
	PIN pin_895
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.429282868525675 0 56.679282868525675 0.25 ;
		END PORT
	END pin_895
	PIN pin_896
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.74900398406352 0 56.99900398406352 0.25 ;
		END PORT
	END pin_896
	PIN pin_897
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.068725099601366 0 57.318725099601366 0.25 ;
		END PORT
	END pin_897
	PIN pin_898
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.38844621513921 0 57.63844621513921 0.25 ;
		END PORT
	END pin_898
	PIN pin_899
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.70816733067706 0 57.95816733067706 0.25 ;
		END PORT
	END pin_899
	PIN pin_900
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.0278884462149 0 58.2778884462149 0.25 ;
		END PORT
	END pin_900
	PIN pin_901
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.34760956175275 0 58.59760956175275 0.25 ;
		END PORT
	END pin_901
	PIN pin_902
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.66733067729059 0 58.91733067729059 0.25 ;
		END PORT
	END pin_902
	PIN pin_903
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.98705179282844 0 59.23705179282844 0.25 ;
		END PORT
	END pin_903
	PIN pin_904
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 59.306772908366284 0 59.556772908366284 0.25 ;
		END PORT
	END pin_904
	PIN pin_905
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 59.62649402390413 0 59.87649402390413 0.25 ;
		END PORT
	END pin_905
	PIN pin_906
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 59.946215139441975 0 60.196215139441975 0.25 ;
		END PORT
	END pin_906
	PIN pin_907
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.26593625497982 0 60.51593625497982 0.25 ;
		END PORT
	END pin_907
	PIN pin_908
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.585657370517666 0 60.835657370517666 0.25 ;
		END PORT
	END pin_908
	PIN pin_909
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 60.90537848605551 0 61.15537848605551 0.25 ;
		END PORT
	END pin_909
	PIN pin_910
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 61.22509960159336 0 61.47509960159336 0.25 ;
		END PORT
	END pin_910
	PIN pin_911
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 61.5448207171312 0 61.7948207171312 0.25 ;
		END PORT
	END pin_911
	PIN pin_912
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 61.86454183266905 0 62.11454183266905 0.25 ;
		END PORT
	END pin_912
	PIN pin_913
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 62.18426294820689 0 62.43426294820689 0.25 ;
		END PORT
	END pin_913
	PIN pin_914
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.50398406374474 0 62.75398406374474 0.25 ;
		END PORT
	END pin_914
	PIN pin_915
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 62.823705179282584 0 63.073705179282584 0.25 ;
		END PORT
	END pin_915
	PIN pin_916
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.14342629482043 0 63.39342629482043 0.25 ;
		END PORT
	END pin_916
	PIN pin_917
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 63.463147410358275 0 63.713147410358275 0.25 ;
		END PORT
	END pin_917
	PIN pin_918
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 63.78286852589612 0 64.03286852589612 0.25 ;
		END PORT
	END pin_918
	PIN pin_919
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 64.10258964143397 0 64.35258964143397 0.25 ;
		END PORT
	END pin_919
	PIN pin_920
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 64.42231075697181 0 64.67231075697181 0.25 ;
		END PORT
	END pin_920
	PIN pin_921
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.74203187250966 0 64.99203187250966 0.25 ;
		END PORT
	END pin_921
	PIN pin_922
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 65.0617529880475 0 65.3117529880475 0.25 ;
		END PORT
	END pin_922
	PIN pin_923
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 65.38147410358535 0 65.63147410358535 0.25 ;
		END PORT
	END pin_923
	PIN pin_924
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 65.70119521912319 0 65.95119521912319 0.25 ;
		END PORT
	END pin_924
	PIN pin_925
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.02091633466104 0 66.27091633466104 0.25 ;
		END PORT
	END pin_925
	PIN pin_926
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.34063745019888 0 66.59063745019888 0.25 ;
		END PORT
	END pin_926
	PIN pin_927
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 66.66035856573673 0 66.91035856573673 0.25 ;
		END PORT
	END pin_927
	PIN pin_928
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.98007968127457 0 67.23007968127457 0.25 ;
		END PORT
	END pin_928
	PIN pin_929
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.29980079681242 0 67.54980079681242 0.25 ;
		END PORT
	END pin_929
	PIN pin_930
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.61952191235027 0 67.86952191235027 0.25 ;
		END PORT
	END pin_930
	PIN pin_931
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.93924302788811 0 68.18924302788811 0.25 ;
		END PORT
	END pin_931
	PIN pin_932
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.25896414342596 0 68.50896414342596 0.25 ;
		END PORT
	END pin_932
	PIN pin_933
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.5786852589638 0 68.8286852589638 0.25 ;
		END PORT
	END pin_933
	PIN pin_934
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 68.89840637450165 0 69.14840637450165 0.25 ;
		END PORT
	END pin_934
	PIN pin_935
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 69.21812749003949 0 69.46812749003949 0.25 ;
		END PORT
	END pin_935
	PIN pin_936
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 69.53784860557734 0 69.78784860557734 0.25 ;
		END PORT
	END pin_936
	PIN pin_937
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 69.85756972111518 0 70.10756972111518 0.25 ;
		END PORT
	END pin_937
	PIN pin_938
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.17729083665303 0 70.42729083665303 0.25 ;
		END PORT
	END pin_938
	PIN pin_939
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 70.49701195219087 0 70.74701195219087 0.25 ;
		END PORT
	END pin_939
	PIN pin_940
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.81673306772872 0 71.06673306772872 0.25 ;
		END PORT
	END pin_940
	PIN pin_941
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 71.13645418326657 0 71.38645418326657 0.25 ;
		END PORT
	END pin_941
	PIN pin_942
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 71.45617529880441 0 71.70617529880441 0.25 ;
		END PORT
	END pin_942
	PIN pin_943
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 71.77589641434226 0 72.02589641434226 0.25 ;
		END PORT
	END pin_943
	PIN pin_944
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 72.0956175298801 0 72.3456175298801 0.25 ;
		END PORT
	END pin_944
	PIN pin_945
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 72.41533864541795 0 72.66533864541795 0.25 ;
		END PORT
	END pin_945
	PIN pin_946
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 72.73505976095579 0 72.98505976095579 0.25 ;
		END PORT
	END pin_946
	PIN pin_947
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.05478087649364 0 73.30478087649364 0.25 ;
		END PORT
	END pin_947
	PIN pin_948
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.37450199203148 0 73.62450199203148 0.25 ;
		END PORT
	END pin_948
	PIN pin_949
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.69422310756933 0 73.94422310756933 0.25 ;
		END PORT
	END pin_949
	PIN pin_950
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.01394422310717 0 74.26394422310717 0.25 ;
		END PORT
	END pin_950
	PIN pin_951
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.33366533864502 0 74.58366533864502 0.25 ;
		END PORT
	END pin_951
	PIN pin_952
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.65338645418286 0 74.90338645418286 0.25 ;
		END PORT
	END pin_952
	PIN pin_953
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 74.97310756972071 0 75.22310756972071 0.25 ;
		END PORT
	END pin_953
	PIN pin_954
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.29282868525856 0 75.54282868525856 0.25 ;
		END PORT
	END pin_954
	PIN pin_955
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 75.6125498007964 0 75.8625498007964 0.25 ;
		END PORT
	END pin_955
	PIN pin_956
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.93227091633425 0 76.18227091633425 0.25 ;
		END PORT
	END pin_956
	PIN pin_957
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.25199203187209 0 76.50199203187209 0.25 ;
		END PORT
	END pin_957
	PIN pin_958
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.57171314740994 0 76.82171314740994 0.25 ;
		END PORT
	END pin_958
	PIN pin_959
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 76.89143426294778 0 77.14143426294778 0.25 ;
		END PORT
	END pin_959
	PIN pin_960
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 77.21115537848563 0 77.46115537848563 0.25 ;
		END PORT
	END pin_960
	PIN pin_961
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.53087649402347 0 77.78087649402347 0.25 ;
		END PORT
	END pin_961
	PIN pin_962
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 77.85059760956132 0 78.10059760956132 0.25 ;
		END PORT
	END pin_962
	PIN pin_963
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 78.17031872509916 0 78.42031872509916 0.25 ;
		END PORT
	END pin_963
	PIN pin_964
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 78.49003984063701 0 78.74003984063701 0.25 ;
		END PORT
	END pin_964
	PIN pin_965
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 78.80976095617486 0 79.05976095617486 0.25 ;
		END PORT
	END pin_965
	PIN pin_966
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.1294820717127 0 79.3794820717127 0.25 ;
		END PORT
	END pin_966
	PIN pin_967
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.44920318725055 0 79.69920318725055 0.25 ;
		END PORT
	END pin_967
	PIN pin_968
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.76892430278839 0 80.01892430278839 0.25 ;
		END PORT
	END pin_968
	PIN pin_969
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 80.08864541832624 0 80.33864541832624 0.25 ;
		END PORT
	END pin_969
	PIN pin_970
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 80.40836653386408 0 80.65836653386408 0.25 ;
		END PORT
	END pin_970
	PIN pin_971
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 80.72808764940193 0 80.97808764940193 0.25 ;
		END PORT
	END pin_971
	PIN pin_972
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 81.04780876493977 0 81.29780876493977 0.25 ;
		END PORT
	END pin_972
	PIN pin_973
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 81.36752988047762 0 81.61752988047762 0.25 ;
		END PORT
	END pin_973
	PIN pin_974
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 81.68725099601546 0 81.93725099601546 0.25 ;
		END PORT
	END pin_974
	PIN pin_975
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.00697211155331 0 82.25697211155331 0.25 ;
		END PORT
	END pin_975
	PIN pin_976
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.32669322709116 0 82.57669322709116 0.25 ;
		END PORT
	END pin_976
	PIN pin_977
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.646414342629 0 82.896414342629 0.25 ;
		END PORT
	END pin_977
	PIN pin_978
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.96613545816685 0 83.21613545816685 0.25 ;
		END PORT
	END pin_978
	PIN pin_979
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 83.28585657370469 0 83.53585657370469 0.25 ;
		END PORT
	END pin_979
	PIN pin_980
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.60557768924254 0 83.85557768924254 0.25 ;
		END PORT
	END pin_980
	PIN pin_981
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.92529880478038 0 84.17529880478038 0.25 ;
		END PORT
	END pin_981
	PIN pin_982
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 84.24501992031823 0 84.49501992031823 0.25 ;
		END PORT
	END pin_982
	PIN pin_983
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 84.56474103585607 0 84.81474103585607 0.25 ;
		END PORT
	END pin_983
	PIN pin_984
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 84.88446215139392 0 85.13446215139392 0.25 ;
		END PORT
	END pin_984
	PIN pin_985
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 85.20418326693176 0 85.45418326693176 0.25 ;
		END PORT
	END pin_985
	PIN pin_986
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 85.52390438246961 0 85.77390438246961 0.25 ;
		END PORT
	END pin_986
	PIN pin_987
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 85.84362549800746 0 86.09362549800746 0.25 ;
		END PORT
	END pin_987
	PIN pin_988
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.1633466135453 0 86.4133466135453 0.25 ;
		END PORT
	END pin_988
	PIN pin_989
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.48306772908315 0 86.73306772908315 0.25 ;
		END PORT
	END pin_989
	PIN pin_990
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 86.80278884462099 0 87.05278884462099 0.25 ;
		END PORT
	END pin_990
	PIN pin_991
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.12250996015884 0 87.37250996015884 0.25 ;
		END PORT
	END pin_991
	PIN pin_992
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.44223107569668 0 87.69223107569668 0.25 ;
		END PORT
	END pin_992
	PIN pin_993
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 87.76195219123453 0 88.01195219123453 0.25 ;
		END PORT
	END pin_993
	PIN pin_994
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.08167330677237 0 88.33167330677237 0.25 ;
		END PORT
	END pin_994
	PIN pin_995
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.40139442231022 0 88.65139442231022 0.25 ;
		END PORT
	END pin_995
	PIN pin_996
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.72111553784806 0 88.97111553784806 0.25 ;
		END PORT
	END pin_996
	PIN pin_997
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.04083665338591 0 89.29083665338591 0.25 ;
		END PORT
	END pin_997
	PIN pin_998
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 89.36055776892375 0 89.61055776892375 0.25 ;
		END PORT
	END pin_998
	PIN pin_999
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.6802788844616 0 89.9302788844616 0.25 ;
		END PORT
	END pin_999
END MACRO
MACRO cell_2
	SIZE 100 BY 100 ;
	PIN pin_0
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 89.68027888446215 0.25 89.93027888446215 ;
		END PORT
	END pin_0
	PIN pin_1
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 89.36055776892431 0.25 89.61055776892431 ;
		END PORT
	END pin_1
	PIN pin_2
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 89.04083665338646 0.25 89.29083665338646 ;
		END PORT
	END pin_2
	PIN pin_3
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 88.72111553784862 0.25 88.97111553784862 ;
		END PORT
	END pin_3
	PIN pin_4
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 88.40139442231077 0.25 88.65139442231077 ;
		END PORT
	END pin_4
	PIN pin_5
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 88.08167330677293 0.25 88.33167330677293 ;
		END PORT
	END pin_5
	PIN pin_6
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 87.76195219123508 0.25 88.01195219123508 ;
		END PORT
	END pin_6
	PIN pin_7
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 87.44223107569724 0.25 87.69223107569724 ;
		END PORT
	END pin_7
	PIN pin_8
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 87.12250996015939 0.25 87.37250996015939 ;
		END PORT
	END pin_8
	PIN pin_9
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 86.80278884462155 0.25 87.05278884462155 ;
		END PORT
	END pin_9
	PIN pin_10
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 86.4830677290837 0.25 86.7330677290837 ;
		END PORT
	END pin_10
	PIN pin_11
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 86.16334661354585 0.25 86.41334661354585 ;
		END PORT
	END pin_11
	PIN pin_12
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 85.84362549800801 0.25 86.09362549800801 ;
		END PORT
	END pin_12
	PIN pin_13
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 85.52390438247016 0.25 85.77390438247016 ;
		END PORT
	END pin_13
	PIN pin_14
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 85.20418326693232 0.25 85.45418326693232 ;
		END PORT
	END pin_14
	PIN pin_15
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 84.88446215139447 0.25 85.13446215139447 ;
		END PORT
	END pin_15
	PIN pin_16
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 84.56474103585663 0.25 84.81474103585663 ;
		END PORT
	END pin_16
	PIN pin_17
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 84.24501992031878 0.25 84.49501992031878 ;
		END PORT
	END pin_17
	PIN pin_18
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 83.92529880478094 0.25 84.17529880478094 ;
		END PORT
	END pin_18
	PIN pin_19
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 83.60557768924309 0.25 83.85557768924309 ;
		END PORT
	END pin_19
	PIN pin_20
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 83.28585657370525 0.25 83.53585657370525 ;
		END PORT
	END pin_20
	PIN pin_21
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 82.9661354581674 0.25 83.2161354581674 ;
		END PORT
	END pin_21
	PIN pin_22
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 82.64641434262955 0.25 82.89641434262955 ;
		END PORT
	END pin_22
	PIN pin_23
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 82.32669322709171 0.25 82.57669322709171 ;
		END PORT
	END pin_23
	PIN pin_24
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 82.00697211155386 0.25 82.25697211155386 ;
		END PORT
	END pin_24
	PIN pin_25
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 81.68725099601602 0.25 81.93725099601602 ;
		END PORT
	END pin_25
	PIN pin_26
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 81.36752988047817 0.25 81.61752988047817 ;
		END PORT
	END pin_26
	PIN pin_27
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 81.04780876494033 0.25 81.29780876494033 ;
		END PORT
	END pin_27
	PIN pin_28
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 80.72808764940248 0.25 80.97808764940248 ;
		END PORT
	END pin_28
	PIN pin_29
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 80.40836653386464 0.25 80.65836653386464 ;
		END PORT
	END pin_29
	PIN pin_30
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 80.08864541832679 0.25 80.33864541832679 ;
		END PORT
	END pin_30
	PIN pin_31
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 79.76892430278895 0.25 80.01892430278895 ;
		END PORT
	END pin_31
	PIN pin_32
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 79.4492031872511 0.25 79.6992031872511 ;
		END PORT
	END pin_32
	PIN pin_33
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 79.12948207171326 0.25 79.37948207171326 ;
		END PORT
	END pin_33
	PIN pin_34
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 78.80976095617541 0.25 79.05976095617541 ;
		END PORT
	END pin_34
	PIN pin_35
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 78.49003984063756 0.25 78.74003984063756 ;
		END PORT
	END pin_35
	PIN pin_36
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 78.17031872509972 0.25 78.42031872509972 ;
		END PORT
	END pin_36
	PIN pin_37
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 77.85059760956187 0.25 78.10059760956187 ;
		END PORT
	END pin_37
	PIN pin_38
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 77.53087649402403 0.25 77.78087649402403 ;
		END PORT
	END pin_38
	PIN pin_39
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 77.21115537848618 0.25 77.46115537848618 ;
		END PORT
	END pin_39
	PIN pin_40
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 76.89143426294834 0.25 77.14143426294834 ;
		END PORT
	END pin_40
	PIN pin_41
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 76.57171314741049 0.25 76.82171314741049 ;
		END PORT
	END pin_41
	PIN pin_42
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 76.25199203187265 0.25 76.50199203187265 ;
		END PORT
	END pin_42
	PIN pin_43
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 75.9322709163348 0.25 76.1822709163348 ;
		END PORT
	END pin_43
	PIN pin_44
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 75.61254980079696 0.25 75.86254980079696 ;
		END PORT
	END pin_44
	PIN pin_45
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 75.29282868525911 0.25 75.54282868525911 ;
		END PORT
	END pin_45
	PIN pin_46
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 74.97310756972126 0.25 75.22310756972126 ;
		END PORT
	END pin_46
	PIN pin_47
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 74.65338645418342 0.25 74.90338645418342 ;
		END PORT
	END pin_47
	PIN pin_48
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 74.33366533864557 0.25 74.58366533864557 ;
		END PORT
	END pin_48
	PIN pin_49
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 74.01394422310773 0.25 74.26394422310773 ;
		END PORT
	END pin_49
	PIN pin_50
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 73.69422310756988 0.25 73.94422310756988 ;
		END PORT
	END pin_50
	PIN pin_51
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 73.37450199203204 0.25 73.62450199203204 ;
		END PORT
	END pin_51
	PIN pin_52
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 73.05478087649419 0.25 73.30478087649419 ;
		END PORT
	END pin_52
	PIN pin_53
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 72.73505976095635 0.25 72.98505976095635 ;
		END PORT
	END pin_53
	PIN pin_54
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 72.4153386454185 0.25 72.6653386454185 ;
		END PORT
	END pin_54
	PIN pin_55
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 72.09561752988066 0.25 72.34561752988066 ;
		END PORT
	END pin_55
	PIN pin_56
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 71.77589641434281 0.25 72.02589641434281 ;
		END PORT
	END pin_56
	PIN pin_57
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 71.45617529880496 0.25 71.70617529880496 ;
		END PORT
	END pin_57
	PIN pin_58
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 71.13645418326712 0.25 71.38645418326712 ;
		END PORT
	END pin_58
	PIN pin_59
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 70.81673306772927 0.25 71.06673306772927 ;
		END PORT
	END pin_59
	PIN pin_60
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 70.49701195219143 0.25 70.74701195219143 ;
		END PORT
	END pin_60
	PIN pin_61
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 70.17729083665358 0.25 70.42729083665358 ;
		END PORT
	END pin_61
	PIN pin_62
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 69.85756972111574 0.25 70.10756972111574 ;
		END PORT
	END pin_62
	PIN pin_63
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 69.53784860557789 0.25 69.78784860557789 ;
		END PORT
	END pin_63
	PIN pin_64
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 69.21812749004005 0.25 69.46812749004005 ;
		END PORT
	END pin_64
	PIN pin_65
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 68.8984063745022 0.25 69.1484063745022 ;
		END PORT
	END pin_65
	PIN pin_66
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 68.57868525896436 0.25 68.82868525896436 ;
		END PORT
	END pin_66
	PIN pin_67
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 68.25896414342651 0.25 68.50896414342651 ;
		END PORT
	END pin_67
	PIN pin_68
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 67.93924302788866 0.25 68.18924302788866 ;
		END PORT
	END pin_68
	PIN pin_69
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 67.61952191235082 0.25 67.86952191235082 ;
		END PORT
	END pin_69
	PIN pin_70
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 67.29980079681297 0.25 67.54980079681297 ;
		END PORT
	END pin_70
	PIN pin_71
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 66.98007968127513 0.25 67.23007968127513 ;
		END PORT
	END pin_71
	PIN pin_72
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 66.66035856573728 0.25 66.91035856573728 ;
		END PORT
	END pin_72
	PIN pin_73
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 66.34063745019944 0.25 66.59063745019944 ;
		END PORT
	END pin_73
	PIN pin_74
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 66.02091633466159 0.25 66.27091633466159 ;
		END PORT
	END pin_74
	PIN pin_75
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 65.70119521912375 0.25 65.95119521912375 ;
		END PORT
	END pin_75
	PIN pin_76
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 65.3814741035859 0.25 65.6314741035859 ;
		END PORT
	END pin_76
	PIN pin_77
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 65.06175298804806 0.25 65.31175298804806 ;
		END PORT
	END pin_77
	PIN pin_78
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 64.74203187251021 0.25 64.99203187251021 ;
		END PORT
	END pin_78
	PIN pin_79
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 64.42231075697237 0.25 64.67231075697237 ;
		END PORT
	END pin_79
	PIN pin_80
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 64.10258964143452 0.25 64.35258964143452 ;
		END PORT
	END pin_80
	PIN pin_81
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 63.782868525896674 0.25 64.03286852589667 ;
		END PORT
	END pin_81
	PIN pin_82
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 63.46314741035883 0.25 63.71314741035883 ;
		END PORT
	END pin_82
	PIN pin_83
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 63.14342629482098 0.25 63.39342629482098 ;
		END PORT
	END pin_83
	PIN pin_84
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 62.82370517928314 0.25 63.07370517928314 ;
		END PORT
	END pin_84
	PIN pin_85
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 62.50398406374529 0.25 62.75398406374529 ;
		END PORT
	END pin_85
	PIN pin_86
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 62.18426294820745 0.25 62.43426294820745 ;
		END PORT
	END pin_86
	PIN pin_87
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 61.8645418326696 0.25 62.1145418326696 ;
		END PORT
	END pin_87
	PIN pin_88
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 61.544820717131756 0.25 61.794820717131756 ;
		END PORT
	END pin_88
	PIN pin_89
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 61.22509960159391 0.25 61.47509960159391 ;
		END PORT
	END pin_89
	PIN pin_90
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 60.905378486056065 0.25 61.155378486056065 ;
		END PORT
	END pin_90
	PIN pin_91
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 60.58565737051822 0.25 60.83565737051822 ;
		END PORT
	END pin_91
	PIN pin_92
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 60.265936254980375 0.25 60.515936254980375 ;
		END PORT
	END pin_92
	PIN pin_93
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 59.94621513944253 0.25 60.19621513944253 ;
		END PORT
	END pin_93
	PIN pin_94
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 59.626494023904684 0.25 59.876494023904684 ;
		END PORT
	END pin_94
	PIN pin_95
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 59.30677290836684 0.25 59.55677290836684 ;
		END PORT
	END pin_95
	PIN pin_96
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.98705179282899 0.25 59.23705179282899 ;
		END PORT
	END pin_96
	PIN pin_97
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 58.66733067729115 0.25 58.91733067729115 ;
		END PORT
	END pin_97
	PIN pin_98
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.3476095617533 0.25 58.5976095617533 ;
		END PORT
	END pin_98
	PIN pin_99
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 58.02788844621546 0.25 58.27788844621546 ;
		END PORT
	END pin_99
	PIN pin_100
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 57.70816733067761 0.25 57.95816733067761 ;
		END PORT
	END pin_100
	PIN pin_101
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 57.388446215139766 0.25 57.638446215139766 ;
		END PORT
	END pin_101
	PIN pin_102
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 57.06872509960192 0.25 57.31872509960192 ;
		END PORT
	END pin_102
	PIN pin_103
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 56.749003984064075 0.25 56.999003984064075 ;
		END PORT
	END pin_103
	PIN pin_104
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 56.42928286852623 0.25 56.67928286852623 ;
		END PORT
	END pin_104
	PIN pin_105
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 56.109561752988384 0.25 56.359561752988384 ;
		END PORT
	END pin_105
	PIN pin_106
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 55.78984063745054 0.25 56.03984063745054 ;
		END PORT
	END pin_106
	PIN pin_107
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 55.47011952191269 0.25 55.72011952191269 ;
		END PORT
	END pin_107
	PIN pin_108
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 55.15039840637485 0.25 55.40039840637485 ;
		END PORT
	END pin_108
	PIN pin_109
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 54.830677290837 0.25 55.080677290837 ;
		END PORT
	END pin_109
	PIN pin_110
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 54.51095617529916 0.25 54.76095617529916 ;
		END PORT
	END pin_110
	PIN pin_111
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 54.19123505976131 0.25 54.44123505976131 ;
		END PORT
	END pin_111
	PIN pin_112
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 53.871513944223466 0.25 54.121513944223466 ;
		END PORT
	END pin_112
	PIN pin_113
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 53.55179282868562 0.25 53.80179282868562 ;
		END PORT
	END pin_113
	PIN pin_114
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 53.232071713147775 0.25 53.482071713147775 ;
		END PORT
	END pin_114
	PIN pin_115
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 52.91235059760993 0.25 53.16235059760993 ;
		END PORT
	END pin_115
	PIN pin_116
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 52.592629482072084 0.25 52.842629482072084 ;
		END PORT
	END pin_116
	PIN pin_117
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 52.27290836653424 0.25 52.52290836653424 ;
		END PORT
	END pin_117
	PIN pin_118
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 51.95318725099639 0.25 52.20318725099639 ;
		END PORT
	END pin_118
	PIN pin_119
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 51.63346613545855 0.25 51.88346613545855 ;
		END PORT
	END pin_119
	PIN pin_120
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 51.3137450199207 0.25 51.5637450199207 ;
		END PORT
	END pin_120
	PIN pin_121
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 50.99402390438286 0.25 51.24402390438286 ;
		END PORT
	END pin_121
	PIN pin_122
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 50.67430278884501 0.25 50.92430278884501 ;
		END PORT
	END pin_122
	PIN pin_123
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 50.354581673307166 0.25 50.604581673307166 ;
		END PORT
	END pin_123
	PIN pin_124
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 50.03486055776932 0.25 50.28486055776932 ;
		END PORT
	END pin_124
	PIN pin_125
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 49.715139442231475 0.25 49.965139442231475 ;
		END PORT
	END pin_125
	PIN pin_126
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 49.39541832669363 0.25 49.64541832669363 ;
		END PORT
	END pin_126
	PIN pin_127
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 49.075697211155784 0.25 49.325697211155784 ;
		END PORT
	END pin_127
	PIN pin_128
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 48.75597609561794 0.25 49.00597609561794 ;
		END PORT
	END pin_128
	PIN pin_129
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 48.43625498008009 0.25 48.68625498008009 ;
		END PORT
	END pin_129
	PIN pin_130
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 48.11653386454225 0.25 48.36653386454225 ;
		END PORT
	END pin_130
	PIN pin_131
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 47.7968127490044 0.25 48.0468127490044 ;
		END PORT
	END pin_131
	PIN pin_132
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 47.47709163346656 0.25 47.72709163346656 ;
		END PORT
	END pin_132
	PIN pin_133
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 47.15737051792871 0.25 47.40737051792871 ;
		END PORT
	END pin_133
	PIN pin_134
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 46.837649402390866 0.25 47.087649402390866 ;
		END PORT
	END pin_134
	PIN pin_135
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 46.51792828685302 0.25 46.76792828685302 ;
		END PORT
	END pin_135
	PIN pin_136
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 46.198207171315175 0.25 46.448207171315175 ;
		END PORT
	END pin_136
	PIN pin_137
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 45.87848605577733 0.25 46.12848605577733 ;
		END PORT
	END pin_137
	PIN pin_138
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 45.558764940239485 0.25 45.808764940239485 ;
		END PORT
	END pin_138
	PIN pin_139
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 45.23904382470164 0.25 45.48904382470164 ;
		END PORT
	END pin_139
	PIN pin_140
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 44.919322709163794 0.25 45.169322709163794 ;
		END PORT
	END pin_140
	PIN pin_141
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 44.59960159362595 0.25 44.84960159362595 ;
		END PORT
	END pin_141
	PIN pin_142
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 44.2798804780881 0.25 44.5298804780881 ;
		END PORT
	END pin_142
	PIN pin_143
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 43.96015936255026 0.25 44.21015936255026 ;
		END PORT
	END pin_143
	PIN pin_144
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 43.64043824701241 0.25 43.89043824701241 ;
		END PORT
	END pin_144
	PIN pin_145
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 43.32071713147457 0.25 43.57071713147457 ;
		END PORT
	END pin_145
	PIN pin_146
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 43.00099601593672 0.25 43.25099601593672 ;
		END PORT
	END pin_146
	PIN pin_147
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 42.681274900398876 0.25 42.931274900398876 ;
		END PORT
	END pin_147
	PIN pin_148
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 42.36155378486103 0.25 42.61155378486103 ;
		END PORT
	END pin_148
	PIN pin_149
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 42.041832669323185 0.25 42.291832669323185 ;
		END PORT
	END pin_149
	PIN pin_150
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 41.72211155378534 0.25 41.97211155378534 ;
		END PORT
	END pin_150
	PIN pin_151
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 41.402390438247494 0.25 41.652390438247494 ;
		END PORT
	END pin_151
	PIN pin_152
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 41.08266932270965 0.25 41.33266932270965 ;
		END PORT
	END pin_152
	PIN pin_153
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 40.7629482071718 0.25 41.0129482071718 ;
		END PORT
	END pin_153
	PIN pin_154
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 40.44322709163396 0.25 40.69322709163396 ;
		END PORT
	END pin_154
	PIN pin_155
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 40.12350597609611 0.25 40.37350597609611 ;
		END PORT
	END pin_155
	PIN pin_156
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 39.80378486055827 0.25 40.05378486055827 ;
		END PORT
	END pin_156
	PIN pin_157
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 39.48406374502042 0.25 39.73406374502042 ;
		END PORT
	END pin_157
	PIN pin_158
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 39.164342629482576 0.25 39.414342629482576 ;
		END PORT
	END pin_158
	PIN pin_159
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 38.84462151394473 0.25 39.09462151394473 ;
		END PORT
	END pin_159
	PIN pin_160
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 38.524900398406885 0.25 38.774900398406885 ;
		END PORT
	END pin_160
	PIN pin_161
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 38.20517928286904 0.25 38.45517928286904 ;
		END PORT
	END pin_161
	PIN pin_162
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 37.885458167331194 0.25 38.135458167331194 ;
		END PORT
	END pin_162
	PIN pin_163
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 37.56573705179335 0.25 37.81573705179335 ;
		END PORT
	END pin_163
	PIN pin_164
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 37.2460159362555 0.25 37.4960159362555 ;
		END PORT
	END pin_164
	PIN pin_165
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 36.92629482071766 0.25 37.17629482071766 ;
		END PORT
	END pin_165
	PIN pin_166
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 36.60657370517981 0.25 36.85657370517981 ;
		END PORT
	END pin_166
	PIN pin_167
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 36.28685258964197 0.25 36.53685258964197 ;
		END PORT
	END pin_167
	PIN pin_168
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 35.96713147410412 0.25 36.21713147410412 ;
		END PORT
	END pin_168
	PIN pin_169
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 35.647410358566276 0.25 35.897410358566276 ;
		END PORT
	END pin_169
	PIN pin_170
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 35.32768924302843 0.25 35.57768924302843 ;
		END PORT
	END pin_170
	PIN pin_171
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 35.007968127490585 0.25 35.257968127490585 ;
		END PORT
	END pin_171
	PIN pin_172
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 34.68824701195274 0.25 34.93824701195274 ;
		END PORT
	END pin_172
	PIN pin_173
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 34.368525896414894 0.25 34.618525896414894 ;
		END PORT
	END pin_173
	PIN pin_174
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 34.04880478087705 0.25 34.29880478087705 ;
		END PORT
	END pin_174
	PIN pin_175
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 33.7290836653392 0.25 33.9790836653392 ;
		END PORT
	END pin_175
	PIN pin_176
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 33.40936254980136 0.25 33.65936254980136 ;
		END PORT
	END pin_176
	PIN pin_177
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 33.08964143426351 0.25 33.33964143426351 ;
		END PORT
	END pin_177
	PIN pin_178
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 32.76992031872567 0.25 33.01992031872567 ;
		END PORT
	END pin_178
	PIN pin_179
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 32.45019920318782 0.25 32.70019920318782 ;
		END PORT
	END pin_179
	PIN pin_180
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 32.130478087649976 0.25 32.380478087649976 ;
		END PORT
	END pin_180
	PIN pin_181
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 31.81075697211213 0.25 32.06075697211213 ;
		END PORT
	END pin_181
	PIN pin_182
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 31.491035856574282 0.25 31.741035856574282 ;
		END PORT
	END pin_182
	PIN pin_183
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 31.171314741036433 0.25 31.421314741036433 ;
		END PORT
	END pin_183
	PIN pin_184
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 30.851593625498584 0.25 31.101593625498584 ;
		END PORT
	END pin_184
	PIN pin_185
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 30.531872509960735 0.25 30.781872509960735 ;
		END PORT
	END pin_185
	PIN pin_186
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 30.212151394422886 0.25 30.462151394422886 ;
		END PORT
	END pin_186
	PIN pin_187
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 29.892430278885037 0.25 30.142430278885037 ;
		END PORT
	END pin_187
	PIN pin_188
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 29.572709163347188 0.25 29.822709163347188 ;
		END PORT
	END pin_188
	PIN pin_189
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 29.25298804780934 0.25 29.50298804780934 ;
		END PORT
	END pin_189
	PIN pin_190
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 28.93326693227149 0.25 29.18326693227149 ;
		END PORT
	END pin_190
	PIN pin_191
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 28.61354581673364 0.25 28.86354581673364 ;
		END PORT
	END pin_191
	PIN pin_192
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 28.293824701195792 0.25 28.543824701195792 ;
		END PORT
	END pin_192
	PIN pin_193
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 27.974103585657943 0.25 28.224103585657943 ;
		END PORT
	END pin_193
	PIN pin_194
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 27.654382470120094 0.25 27.904382470120094 ;
		END PORT
	END pin_194
	PIN pin_195
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 27.334661354582245 0.25 27.584661354582245 ;
		END PORT
	END pin_195
	PIN pin_196
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 27.014940239044396 0.25 27.264940239044396 ;
		END PORT
	END pin_196
	PIN pin_197
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 26.695219123506547 0.25 26.945219123506547 ;
		END PORT
	END pin_197
	PIN pin_198
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 26.375498007968698 0.25 26.625498007968698 ;
		END PORT
	END pin_198
	PIN pin_199
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 26.05577689243085 0.25 26.30577689243085 ;
		END PORT
	END pin_199
	PIN pin_200
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 25.736055776893 0.25 25.986055776893 ;
		END PORT
	END pin_200
	PIN pin_201
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 25.41633466135515 0.25 25.66633466135515 ;
		END PORT
	END pin_201
	PIN pin_202
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 25.096613545817302 0.25 25.346613545817302 ;
		END PORT
	END pin_202
	PIN pin_203
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 24.776892430279453 0.25 25.026892430279453 ;
		END PORT
	END pin_203
	PIN pin_204
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 24.457171314741604 0.25 24.707171314741604 ;
		END PORT
	END pin_204
	PIN pin_205
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 24.137450199203755 0.25 24.387450199203755 ;
		END PORT
	END pin_205
	PIN pin_206
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 23.817729083665906 0.25 24.067729083665906 ;
		END PORT
	END pin_206
	PIN pin_207
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 23.498007968128057 0.25 23.748007968128057 ;
		END PORT
	END pin_207
	PIN pin_208
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 23.178286852590208 0.25 23.428286852590208 ;
		END PORT
	END pin_208
	PIN pin_209
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 22.85856573705236 0.25 23.10856573705236 ;
		END PORT
	END pin_209
	PIN pin_210
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 22.53884462151451 0.25 22.78884462151451 ;
		END PORT
	END pin_210
	PIN pin_211
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 22.21912350597666 0.25 22.46912350597666 ;
		END PORT
	END pin_211
	PIN pin_212
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 21.899402390438812 0.25 22.149402390438812 ;
		END PORT
	END pin_212
	PIN pin_213
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 21.579681274900963 0.25 21.829681274900963 ;
		END PORT
	END pin_213
	PIN pin_214
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 21.259960159363114 0.25 21.509960159363114 ;
		END PORT
	END pin_214
	PIN pin_215
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 20.940239043825265 0.25 21.190239043825265 ;
		END PORT
	END pin_215
	PIN pin_216
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 20.620517928287416 0.25 20.870517928287416 ;
		END PORT
	END pin_216
	PIN pin_217
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 20.300796812749567 0.25 20.550796812749567 ;
		END PORT
	END pin_217
	PIN pin_218
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 19.98107569721172 0.25 20.23107569721172 ;
		END PORT
	END pin_218
	PIN pin_219
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 19.66135458167387 0.25 19.91135458167387 ;
		END PORT
	END pin_219
	PIN pin_220
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 19.34163346613602 0.25 19.59163346613602 ;
		END PORT
	END pin_220
	PIN pin_221
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 19.02191235059817 0.25 19.27191235059817 ;
		END PORT
	END pin_221
	PIN pin_222
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 18.702191235060322 0.25 18.952191235060322 ;
		END PORT
	END pin_222
	PIN pin_223
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 18.382470119522473 0.25 18.632470119522473 ;
		END PORT
	END pin_223
	PIN pin_224
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 18.062749003984624 0.25 18.312749003984624 ;
		END PORT
	END pin_224
	PIN pin_225
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 17.743027888446775 0.25 17.993027888446775 ;
		END PORT
	END pin_225
	PIN pin_226
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 17.423306772908926 0.25 17.673306772908926 ;
		END PORT
	END pin_226
	PIN pin_227
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 17.103585657371077 0.25 17.353585657371077 ;
		END PORT
	END pin_227
	PIN pin_228
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 16.78386454183323 0.25 17.03386454183323 ;
		END PORT
	END pin_228
	PIN pin_229
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 16.46414342629538 0.25 16.71414342629538 ;
		END PORT
	END pin_229
	PIN pin_230
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 16.14442231075753 0.25 16.39442231075753 ;
		END PORT
	END pin_230
	PIN pin_231
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 15.824701195219681 0.25 16.07470119521968 ;
		END PORT
	END pin_231
	PIN pin_232
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 15.504980079681832 0.25 15.754980079681832 ;
		END PORT
	END pin_232
	PIN pin_233
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 15.185258964143983 0.25 15.435258964143983 ;
		END PORT
	END pin_233
	PIN pin_234
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 14.865537848606134 0.25 15.115537848606134 ;
		END PORT
	END pin_234
	PIN pin_235
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 14.545816733068285 0.25 14.795816733068285 ;
		END PORT
	END pin_235
	PIN pin_236
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 14.226095617530436 0.25 14.476095617530436 ;
		END PORT
	END pin_236
	PIN pin_237
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 13.906374501992588 0.25 14.156374501992588 ;
		END PORT
	END pin_237
	PIN pin_238
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 13.586653386454739 0.25 13.836653386454739 ;
		END PORT
	END pin_238
	PIN pin_239
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 13.26693227091689 0.25 13.51693227091689 ;
		END PORT
	END pin_239
	PIN pin_240
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 12.94721115537904 0.25 13.19721115537904 ;
		END PORT
	END pin_240
	PIN pin_241
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 12.627490039841192 0.25 12.877490039841192 ;
		END PORT
	END pin_241
	PIN pin_242
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 12.307768924303343 0.25 12.557768924303343 ;
		END PORT
	END pin_242
	PIN pin_243
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 11.988047808765494 0.25 12.238047808765494 ;
		END PORT
	END pin_243
	PIN pin_244
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 11.668326693227645 0.25 11.918326693227645 ;
		END PORT
	END pin_244
	PIN pin_245
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 11.348605577689796 0.25 11.598605577689796 ;
		END PORT
	END pin_245
	PIN pin_246
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 11.028884462151947 0.25 11.278884462151947 ;
		END PORT
	END pin_246
	PIN pin_247
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 10.709163346614098 0.25 10.959163346614098 ;
		END PORT
	END pin_247
	PIN pin_248
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 0 10.389442231076249 0.25 10.639442231076249 ;
		END PORT
	END pin_248
	PIN pin_249
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 10.0697211155384 0.25 10.3197211155384 ;
		END PORT
	END pin_249
	PIN pin_250
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.069721115537849 100 10.319721115537849 ;
		END PORT
	END pin_250
	PIN pin_251
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.389442231075698 100 10.639442231075698 ;
		END PORT
	END pin_251
	PIN pin_252
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 10.709163346613547 100 10.959163346613547 ;
		END PORT
	END pin_252
	PIN pin_253
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.028884462151396 100 11.278884462151396 ;
		END PORT
	END pin_253
	PIN pin_254
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.348605577689245 100 11.598605577689245 ;
		END PORT
	END pin_254
	PIN pin_255
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.668326693227094 100 11.918326693227094 ;
		END PORT
	END pin_255
	PIN pin_256
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 11.988047808764943 100 12.238047808764943 ;
		END PORT
	END pin_256
	PIN pin_257
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.307768924302792 100 12.557768924302792 ;
		END PORT
	END pin_257
	PIN pin_258
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.627490039840641 100 12.877490039840641 ;
		END PORT
	END pin_258
	PIN pin_259
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 12.94721115537849 100 13.19721115537849 ;
		END PORT
	END pin_259
	PIN pin_260
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.266932270916339 100 13.516932270916339 ;
		END PORT
	END pin_260
	PIN pin_261
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.586653386454188 100 13.836653386454188 ;
		END PORT
	END pin_261
	PIN pin_262
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 13.906374501992037 100 14.156374501992037 ;
		END PORT
	END pin_262
	PIN pin_263
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.226095617529886 100 14.476095617529886 ;
		END PORT
	END pin_263
	PIN pin_264
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.545816733067735 100 14.795816733067735 ;
		END PORT
	END pin_264
	PIN pin_265
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 14.865537848605584 100 15.115537848605584 ;
		END PORT
	END pin_265
	PIN pin_266
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.185258964143433 100 15.435258964143433 ;
		END PORT
	END pin_266
	PIN pin_267
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.504980079681282 100 15.754980079681282 ;
		END PORT
	END pin_267
	PIN pin_268
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 15.82470119521913 100 16.07470119521913 ;
		END PORT
	END pin_268
	PIN pin_269
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.14442231075698 100 16.39442231075698 ;
		END PORT
	END pin_269
	PIN pin_270
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.46414342629483 100 16.71414342629483 ;
		END PORT
	END pin_270
	PIN pin_271
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 16.783864541832678 100 17.033864541832678 ;
		END PORT
	END pin_271
	PIN pin_272
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.103585657370527 100 17.353585657370527 ;
		END PORT
	END pin_272
	PIN pin_273
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.423306772908376 100 17.673306772908376 ;
		END PORT
	END pin_273
	PIN pin_274
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 17.743027888446225 100 17.993027888446225 ;
		END PORT
	END pin_274
	PIN pin_275
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.062749003984074 100 18.312749003984074 ;
		END PORT
	END pin_275
	PIN pin_276
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.382470119521923 100 18.632470119521923 ;
		END PORT
	END pin_276
	PIN pin_277
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 18.70219123505977 100 18.95219123505977 ;
		END PORT
	END pin_277
	PIN pin_278
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.02191235059762 100 19.27191235059762 ;
		END PORT
	END pin_278
	PIN pin_279
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.34163346613547 100 19.59163346613547 ;
		END PORT
	END pin_279
	PIN pin_280
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.66135458167332 100 19.91135458167332 ;
		END PORT
	END pin_280
	PIN pin_281
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 19.981075697211168 100 20.231075697211168 ;
		END PORT
	END pin_281
	PIN pin_282
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.300796812749017 100 20.550796812749017 ;
		END PORT
	END pin_282
	PIN pin_283
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.620517928286866 100 20.870517928286866 ;
		END PORT
	END pin_283
	PIN pin_284
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 20.940239043824715 100 21.190239043824715 ;
		END PORT
	END pin_284
	PIN pin_285
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.259960159362564 100 21.509960159362564 ;
		END PORT
	END pin_285
	PIN pin_286
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.579681274900413 100 21.829681274900413 ;
		END PORT
	END pin_286
	PIN pin_287
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 21.89940239043826 100 22.14940239043826 ;
		END PORT
	END pin_287
	PIN pin_288
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.21912350597611 100 22.46912350597611 ;
		END PORT
	END pin_288
	PIN pin_289
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.53884462151396 100 22.78884462151396 ;
		END PORT
	END pin_289
	PIN pin_290
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 22.85856573705181 100 23.10856573705181 ;
		END PORT
	END pin_290
	PIN pin_291
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.178286852589657 100 23.428286852589657 ;
		END PORT
	END pin_291
	PIN pin_292
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.498007968127506 100 23.748007968127506 ;
		END PORT
	END pin_292
	PIN pin_293
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 23.817729083665355 100 24.067729083665355 ;
		END PORT
	END pin_293
	PIN pin_294
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.137450199203204 100 24.387450199203204 ;
		END PORT
	END pin_294
	PIN pin_295
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.457171314741053 100 24.707171314741053 ;
		END PORT
	END pin_295
	PIN pin_296
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 24.776892430278902 100 25.026892430278902 ;
		END PORT
	END pin_296
	PIN pin_297
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.09661354581675 100 25.34661354581675 ;
		END PORT
	END pin_297
	PIN pin_298
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.4163346613546 100 25.6663346613546 ;
		END PORT
	END pin_298
	PIN pin_299
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 25.73605577689245 100 25.98605577689245 ;
		END PORT
	END pin_299
	PIN pin_300
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.0557768924303 100 26.3057768924303 ;
		END PORT
	END pin_300
	PIN pin_301
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.375498007968147 100 26.625498007968147 ;
		END PORT
	END pin_301
	PIN pin_302
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 26.695219123505996 100 26.945219123505996 ;
		END PORT
	END pin_302
	PIN pin_303
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.014940239043845 100 27.264940239043845 ;
		END PORT
	END pin_303
	PIN pin_304
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.334661354581694 100 27.584661354581694 ;
		END PORT
	END pin_304
	PIN pin_305
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.654382470119543 100 27.904382470119543 ;
		END PORT
	END pin_305
	PIN pin_306
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 27.974103585657392 100 28.224103585657392 ;
		END PORT
	END pin_306
	PIN pin_307
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.29382470119524 100 28.54382470119524 ;
		END PORT
	END pin_307
	PIN pin_308
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.61354581673309 100 28.86354581673309 ;
		END PORT
	END pin_308
	PIN pin_309
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 28.93326693227094 100 29.18326693227094 ;
		END PORT
	END pin_309
	PIN pin_310
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.25298804780879 100 29.50298804780879 ;
		END PORT
	END pin_310
	PIN pin_311
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.572709163346637 100 29.822709163346637 ;
		END PORT
	END pin_311
	PIN pin_312
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 29.892430278884486 100 30.142430278884486 ;
		END PORT
	END pin_312
	PIN pin_313
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.212151394422335 100 30.462151394422335 ;
		END PORT
	END pin_313
	PIN pin_314
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.531872509960184 100 30.781872509960184 ;
		END PORT
	END pin_314
	PIN pin_315
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 30.851593625498033 100 31.101593625498033 ;
		END PORT
	END pin_315
	PIN pin_316
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.171314741035882 100 31.421314741035882 ;
		END PORT
	END pin_316
	PIN pin_317
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.49103585657373 100 31.74103585657373 ;
		END PORT
	END pin_317
	PIN pin_318
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 31.81075697211158 100 32.06075697211158 ;
		END PORT
	END pin_318
	PIN pin_319
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.13047808764942 100 32.38047808764942 ;
		END PORT
	END pin_319
	PIN pin_320
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.45019920318727 100 32.70019920318727 ;
		END PORT
	END pin_320
	PIN pin_321
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 32.76992031872511 100 33.01992031872511 ;
		END PORT
	END pin_321
	PIN pin_322
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.08964143426296 100 33.33964143426296 ;
		END PORT
	END pin_322
	PIN pin_323
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.409362549800804 100 33.659362549800804 ;
		END PORT
	END pin_323
	PIN pin_324
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 33.72908366533865 100 33.97908366533865 ;
		END PORT
	END pin_324
	PIN pin_325
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.048804780876495 100 34.298804780876495 ;
		END PORT
	END pin_325
	PIN pin_326
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.36852589641434 100 34.61852589641434 ;
		END PORT
	END pin_326
	PIN pin_327
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 34.688247011952186 100 34.938247011952186 ;
		END PORT
	END pin_327
	PIN pin_328
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.00796812749003 100 35.25796812749003 ;
		END PORT
	END pin_328
	PIN pin_329
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.327689243027876 100 35.577689243027876 ;
		END PORT
	END pin_329
	PIN pin_330
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.64741035856572 100 35.89741035856572 ;
		END PORT
	END pin_330
	PIN pin_331
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 35.96713147410357 100 36.21713147410357 ;
		END PORT
	END pin_331
	PIN pin_332
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.28685258964141 100 36.53685258964141 ;
		END PORT
	END pin_332
	PIN pin_333
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.60657370517926 100 36.85657370517926 ;
		END PORT
	END pin_333
	PIN pin_334
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 36.926294820717104 100 37.176294820717104 ;
		END PORT
	END pin_334
	PIN pin_335
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.24601593625495 100 37.49601593625495 ;
		END PORT
	END pin_335
	PIN pin_336
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.565737051792794 100 37.815737051792794 ;
		END PORT
	END pin_336
	PIN pin_337
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 37.88545816733064 100 38.13545816733064 ;
		END PORT
	END pin_337
	PIN pin_338
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.205179282868485 100 38.455179282868485 ;
		END PORT
	END pin_338
	PIN pin_339
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.52490039840633 100 38.77490039840633 ;
		END PORT
	END pin_339
	PIN pin_340
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 38.844621513944176 100 39.094621513944176 ;
		END PORT
	END pin_340
	PIN pin_341
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.16434262948202 100 39.41434262948202 ;
		END PORT
	END pin_341
	PIN pin_342
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.48406374501987 100 39.73406374501987 ;
		END PORT
	END pin_342
	PIN pin_343
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 39.80378486055771 100 40.05378486055771 ;
		END PORT
	END pin_343
	PIN pin_344
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.12350597609556 100 40.37350597609556 ;
		END PORT
	END pin_344
	PIN pin_345
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.4432270916334 100 40.6932270916334 ;
		END PORT
	END pin_345
	PIN pin_346
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 40.76294820717125 100 41.01294820717125 ;
		END PORT
	END pin_346
	PIN pin_347
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.082669322709094 100 41.332669322709094 ;
		END PORT
	END pin_347
	PIN pin_348
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.40239043824694 100 41.65239043824694 ;
		END PORT
	END pin_348
	PIN pin_349
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 41.722111553784785 100 41.972111553784785 ;
		END PORT
	END pin_349
	PIN pin_350
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.04183266932263 100 42.29183266932263 ;
		END PORT
	END pin_350
	PIN pin_351
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.361553784860476 100 42.611553784860476 ;
		END PORT
	END pin_351
	PIN pin_352
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 42.68127490039832 100 42.93127490039832 ;
		END PORT
	END pin_352
	PIN pin_353
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.00099601593617 100 43.25099601593617 ;
		END PORT
	END pin_353
	PIN pin_354
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.32071713147401 100 43.57071713147401 ;
		END PORT
	END pin_354
	PIN pin_355
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.64043824701186 100 43.89043824701186 ;
		END PORT
	END pin_355
	PIN pin_356
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 43.9601593625497 100 44.2101593625497 ;
		END PORT
	END pin_356
	PIN pin_357
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.27988047808755 100 44.52988047808755 ;
		END PORT
	END pin_357
	PIN pin_358
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.599601593625394 100 44.849601593625394 ;
		END PORT
	END pin_358
	PIN pin_359
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 44.91932270916324 100 45.16932270916324 ;
		END PORT
	END pin_359
	PIN pin_360
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.239043824701085 100 45.489043824701085 ;
		END PORT
	END pin_360
	PIN pin_361
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.55876494023893 100 45.80876494023893 ;
		END PORT
	END pin_361
	PIN pin_362
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 45.878486055776776 100 46.128486055776776 ;
		END PORT
	END pin_362
	PIN pin_363
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.19820717131462 100 46.44820717131462 ;
		END PORT
	END pin_363
	PIN pin_364
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.51792828685247 100 46.76792828685247 ;
		END PORT
	END pin_364
	PIN pin_365
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 46.83764940239031 100 47.08764940239031 ;
		END PORT
	END pin_365
	PIN pin_366
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.15737051792816 100 47.40737051792816 ;
		END PORT
	END pin_366
	PIN pin_367
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.477091633466 100 47.727091633466 ;
		END PORT
	END pin_367
	PIN pin_368
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 47.79681274900385 100 48.04681274900385 ;
		END PORT
	END pin_368
	PIN pin_369
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.116533864541694 100 48.366533864541694 ;
		END PORT
	END pin_369
	PIN pin_370
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.43625498007954 100 48.68625498007954 ;
		END PORT
	END pin_370
	PIN pin_371
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 48.755976095617385 100 49.005976095617385 ;
		END PORT
	END pin_371
	PIN pin_372
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.07569721115523 100 49.32569721115523 ;
		END PORT
	END pin_372
	PIN pin_373
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.395418326693076 100 49.645418326693076 ;
		END PORT
	END pin_373
	PIN pin_374
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 49.71513944223092 100 49.96513944223092 ;
		END PORT
	END pin_374
	PIN pin_375
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.034860557768766 100 50.284860557768766 ;
		END PORT
	END pin_375
	PIN pin_376
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.35458167330661 100 50.60458167330661 ;
		END PORT
	END pin_376
	PIN pin_377
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.67430278884446 100 50.92430278884446 ;
		END PORT
	END pin_377
	PIN pin_378
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 50.9940239043823 100 51.2440239043823 ;
		END PORT
	END pin_378
	PIN pin_379
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.31374501992015 100 51.56374501992015 ;
		END PORT
	END pin_379
	PIN pin_380
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.633466135457994 100 51.883466135457994 ;
		END PORT
	END pin_380
	PIN pin_381
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 51.95318725099584 100 52.20318725099584 ;
		END PORT
	END pin_381
	PIN pin_382
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.272908366533684 100 52.522908366533684 ;
		END PORT
	END pin_382
	PIN pin_383
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.59262948207153 100 52.84262948207153 ;
		END PORT
	END pin_383
	PIN pin_384
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 52.912350597609375 100 53.162350597609375 ;
		END PORT
	END pin_384
	PIN pin_385
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.23207171314722 100 53.48207171314722 ;
		END PORT
	END pin_385
	PIN pin_386
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.551792828685066 100 53.801792828685066 ;
		END PORT
	END pin_386
	PIN pin_387
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 53.87151394422291 100 54.12151394422291 ;
		END PORT
	END pin_387
	PIN pin_388
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.19123505976076 100 54.44123505976076 ;
		END PORT
	END pin_388
	PIN pin_389
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.5109561752986 100 54.7609561752986 ;
		END PORT
	END pin_389
	PIN pin_390
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 54.83067729083645 100 55.08067729083645 ;
		END PORT
	END pin_390
	PIN pin_391
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.15039840637429 100 55.40039840637429 ;
		END PORT
	END pin_391
	PIN pin_392
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.47011952191214 100 55.72011952191214 ;
		END PORT
	END pin_392
	PIN pin_393
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 55.789840637449984 100 56.039840637449984 ;
		END PORT
	END pin_393
	PIN pin_394
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.10956175298783 100 56.35956175298783 ;
		END PORT
	END pin_394
	PIN pin_395
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.429282868525675 100 56.679282868525675 ;
		END PORT
	END pin_395
	PIN pin_396
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 56.74900398406352 100 56.99900398406352 ;
		END PORT
	END pin_396
	PIN pin_397
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.068725099601366 100 57.318725099601366 ;
		END PORT
	END pin_397
	PIN pin_398
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.38844621513921 100 57.63844621513921 ;
		END PORT
	END pin_398
	PIN pin_399
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 57.70816733067706 100 57.95816733067706 ;
		END PORT
	END pin_399
	PIN pin_400
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.0278884462149 100 58.2778884462149 ;
		END PORT
	END pin_400
	PIN pin_401
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.34760956175275 100 58.59760956175275 ;
		END PORT
	END pin_401
	PIN pin_402
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.66733067729059 100 58.91733067729059 ;
		END PORT
	END pin_402
	PIN pin_403
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 58.98705179282844 100 59.23705179282844 ;
		END PORT
	END pin_403
	PIN pin_404
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.306772908366284 100 59.556772908366284 ;
		END PORT
	END pin_404
	PIN pin_405
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.62649402390413 100 59.87649402390413 ;
		END PORT
	END pin_405
	PIN pin_406
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 59.946215139441975 100 60.196215139441975 ;
		END PORT
	END pin_406
	PIN pin_407
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.26593625497982 100 60.51593625497982 ;
		END PORT
	END pin_407
	PIN pin_408
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.585657370517666 100 60.835657370517666 ;
		END PORT
	END pin_408
	PIN pin_409
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 60.90537848605551 100 61.15537848605551 ;
		END PORT
	END pin_409
	PIN pin_410
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.22509960159336 100 61.47509960159336 ;
		END PORT
	END pin_410
	PIN pin_411
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.5448207171312 100 61.7948207171312 ;
		END PORT
	END pin_411
	PIN pin_412
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 61.86454183266905 100 62.11454183266905 ;
		END PORT
	END pin_412
	PIN pin_413
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.18426294820689 100 62.43426294820689 ;
		END PORT
	END pin_413
	PIN pin_414
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.50398406374474 100 62.75398406374474 ;
		END PORT
	END pin_414
	PIN pin_415
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 62.823705179282584 100 63.073705179282584 ;
		END PORT
	END pin_415
	PIN pin_416
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.14342629482043 100 63.39342629482043 ;
		END PORT
	END pin_416
	PIN pin_417
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.463147410358275 100 63.713147410358275 ;
		END PORT
	END pin_417
	PIN pin_418
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 63.78286852589612 100 64.03286852589612 ;
		END PORT
	END pin_418
	PIN pin_419
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.10258964143397 100 64.35258964143397 ;
		END PORT
	END pin_419
	PIN pin_420
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.42231075697181 100 64.67231075697181 ;
		END PORT
	END pin_420
	PIN pin_421
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 64.74203187250966 100 64.99203187250966 ;
		END PORT
	END pin_421
	PIN pin_422
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.0617529880475 100 65.3117529880475 ;
		END PORT
	END pin_422
	PIN pin_423
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.38147410358535 100 65.63147410358535 ;
		END PORT
	END pin_423
	PIN pin_424
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 65.70119521912319 100 65.95119521912319 ;
		END PORT
	END pin_424
	PIN pin_425
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.02091633466104 100 66.27091633466104 ;
		END PORT
	END pin_425
	PIN pin_426
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.34063745019888 100 66.59063745019888 ;
		END PORT
	END pin_426
	PIN pin_427
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.66035856573673 100 66.91035856573673 ;
		END PORT
	END pin_427
	PIN pin_428
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 66.98007968127457 100 67.23007968127457 ;
		END PORT
	END pin_428
	PIN pin_429
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.29980079681242 100 67.54980079681242 ;
		END PORT
	END pin_429
	PIN pin_430
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.61952191235027 100 67.86952191235027 ;
		END PORT
	END pin_430
	PIN pin_431
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 67.93924302788811 100 68.18924302788811 ;
		END PORT
	END pin_431
	PIN pin_432
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.25896414342596 100 68.50896414342596 ;
		END PORT
	END pin_432
	PIN pin_433
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.5786852589638 100 68.8286852589638 ;
		END PORT
	END pin_433
	PIN pin_434
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 68.89840637450165 100 69.14840637450165 ;
		END PORT
	END pin_434
	PIN pin_435
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.21812749003949 100 69.46812749003949 ;
		END PORT
	END pin_435
	PIN pin_436
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.53784860557734 100 69.78784860557734 ;
		END PORT
	END pin_436
	PIN pin_437
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 69.85756972111518 100 70.10756972111518 ;
		END PORT
	END pin_437
	PIN pin_438
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.17729083665303 100 70.42729083665303 ;
		END PORT
	END pin_438
	PIN pin_439
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.49701195219087 100 70.74701195219087 ;
		END PORT
	END pin_439
	PIN pin_440
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 70.81673306772872 100 71.06673306772872 ;
		END PORT
	END pin_440
	PIN pin_441
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.13645418326657 100 71.38645418326657 ;
		END PORT
	END pin_441
	PIN pin_442
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.45617529880441 100 71.70617529880441 ;
		END PORT
	END pin_442
	PIN pin_443
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 71.77589641434226 100 72.02589641434226 ;
		END PORT
	END pin_443
	PIN pin_444
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.0956175298801 100 72.3456175298801 ;
		END PORT
	END pin_444
	PIN pin_445
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.41533864541795 100 72.66533864541795 ;
		END PORT
	END pin_445
	PIN pin_446
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 72.73505976095579 100 72.98505976095579 ;
		END PORT
	END pin_446
	PIN pin_447
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.05478087649364 100 73.30478087649364 ;
		END PORT
	END pin_447
	PIN pin_448
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.37450199203148 100 73.62450199203148 ;
		END PORT
	END pin_448
	PIN pin_449
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 73.69422310756933 100 73.94422310756933 ;
		END PORT
	END pin_449
	PIN pin_450
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.01394422310717 100 74.26394422310717 ;
		END PORT
	END pin_450
	PIN pin_451
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.33366533864502 100 74.58366533864502 ;
		END PORT
	END pin_451
	PIN pin_452
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.65338645418286 100 74.90338645418286 ;
		END PORT
	END pin_452
	PIN pin_453
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 74.97310756972071 100 75.22310756972071 ;
		END PORT
	END pin_453
	PIN pin_454
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.29282868525856 100 75.54282868525856 ;
		END PORT
	END pin_454
	PIN pin_455
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.6125498007964 100 75.8625498007964 ;
		END PORT
	END pin_455
	PIN pin_456
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 75.93227091633425 100 76.18227091633425 ;
		END PORT
	END pin_456
	PIN pin_457
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.25199203187209 100 76.50199203187209 ;
		END PORT
	END pin_457
	PIN pin_458
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.57171314740994 100 76.82171314740994 ;
		END PORT
	END pin_458
	PIN pin_459
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 76.89143426294778 100 77.14143426294778 ;
		END PORT
	END pin_459
	PIN pin_460
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.21115537848563 100 77.46115537848563 ;
		END PORT
	END pin_460
	PIN pin_461
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.53087649402347 100 77.78087649402347 ;
		END PORT
	END pin_461
	PIN pin_462
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 77.85059760956132 100 78.10059760956132 ;
		END PORT
	END pin_462
	PIN pin_463
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.17031872509916 100 78.42031872509916 ;
		END PORT
	END pin_463
	PIN pin_464
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.49003984063701 100 78.74003984063701 ;
		END PORT
	END pin_464
	PIN pin_465
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 78.80976095617486 100 79.05976095617486 ;
		END PORT
	END pin_465
	PIN pin_466
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.1294820717127 100 79.3794820717127 ;
		END PORT
	END pin_466
	PIN pin_467
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.44920318725055 100 79.69920318725055 ;
		END PORT
	END pin_467
	PIN pin_468
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 79.76892430278839 100 80.01892430278839 ;
		END PORT
	END pin_468
	PIN pin_469
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.08864541832624 100 80.33864541832624 ;
		END PORT
	END pin_469
	PIN pin_470
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.40836653386408 100 80.65836653386408 ;
		END PORT
	END pin_470
	PIN pin_471
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 80.72808764940193 100 80.97808764940193 ;
		END PORT
	END pin_471
	PIN pin_472
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.04780876493977 100 81.29780876493977 ;
		END PORT
	END pin_472
	PIN pin_473
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.36752988047762 100 81.61752988047762 ;
		END PORT
	END pin_473
	PIN pin_474
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 81.68725099601546 100 81.93725099601546 ;
		END PORT
	END pin_474
	PIN pin_475
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.00697211155331 100 82.25697211155331 ;
		END PORT
	END pin_475
	PIN pin_476
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.32669322709116 100 82.57669322709116 ;
		END PORT
	END pin_476
	PIN pin_477
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.646414342629 100 82.896414342629 ;
		END PORT
	END pin_477
	PIN pin_478
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 82.96613545816685 100 83.21613545816685 ;
		END PORT
	END pin_478
	PIN pin_479
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.28585657370469 100 83.53585657370469 ;
		END PORT
	END pin_479
	PIN pin_480
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.60557768924254 100 83.85557768924254 ;
		END PORT
	END pin_480
	PIN pin_481
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 83.92529880478038 100 84.17529880478038 ;
		END PORT
	END pin_481
	PIN pin_482
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.24501992031823 100 84.49501992031823 ;
		END PORT
	END pin_482
	PIN pin_483
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.56474103585607 100 84.81474103585607 ;
		END PORT
	END pin_483
	PIN pin_484
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 84.88446215139392 100 85.13446215139392 ;
		END PORT
	END pin_484
	PIN pin_485
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.20418326693176 100 85.45418326693176 ;
		END PORT
	END pin_485
	PIN pin_486
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.52390438246961 100 85.77390438246961 ;
		END PORT
	END pin_486
	PIN pin_487
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 85.84362549800746 100 86.09362549800746 ;
		END PORT
	END pin_487
	PIN pin_488
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.1633466135453 100 86.4133466135453 ;
		END PORT
	END pin_488
	PIN pin_489
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.48306772908315 100 86.73306772908315 ;
		END PORT
	END pin_489
	PIN pin_490
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 86.80278884462099 100 87.05278884462099 ;
		END PORT
	END pin_490
	PIN pin_491
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.12250996015884 100 87.37250996015884 ;
		END PORT
	END pin_491
	PIN pin_492
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.44223107569668 100 87.69223107569668 ;
		END PORT
	END pin_492
	PIN pin_493
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 87.76195219123453 100 88.01195219123453 ;
		END PORT
	END pin_493
	PIN pin_494
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.08167330677237 100 88.33167330677237 ;
		END PORT
	END pin_494
	PIN pin_495
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.40139442231022 100 88.65139442231022 ;
		END PORT
	END pin_495
	PIN pin_496
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99.75 88.72111553784806 100 88.97111553784806 ;
		END PORT
	END pin_496
	PIN pin_497
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.04083665338591 100 89.29083665338591 ;
		END PORT
	END pin_497
	PIN pin_498
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.36055776892375 100 89.61055776892375 ;
		END PORT
	END pin_498
	PIN pin_499
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99.75 89.6802788844616 100 89.9302788844616 ;
		END PORT
	END pin_499
	PIN pin_500
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 89.68027888446215 99.75 89.93027888446215 100 ;
		END PORT
	END pin_500
	PIN pin_501
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 89.36055776892431 99.75 89.61055776892431 100 ;
		END PORT
	END pin_501
	PIN pin_502
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 89.04083665338646 99.75 89.29083665338646 100 ;
		END PORT
	END pin_502
	PIN pin_503
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 88.72111553784862 99.75 88.97111553784862 100 ;
		END PORT
	END pin_503
	PIN pin_504
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.40139442231077 99.75 88.65139442231077 100 ;
		END PORT
	END pin_504
	PIN pin_505
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 88.08167330677293 99.75 88.33167330677293 100 ;
		END PORT
	END pin_505
	PIN pin_506
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 87.76195219123508 99.75 88.01195219123508 100 ;
		END PORT
	END pin_506
	PIN pin_507
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 87.44223107569724 99.75 87.69223107569724 100 ;
		END PORT
	END pin_507
	PIN pin_508
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 87.12250996015939 99.75 87.37250996015939 100 ;
		END PORT
	END pin_508
	PIN pin_509
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 86.80278884462155 99.75 87.05278884462155 100 ;
		END PORT
	END pin_509
	PIN pin_510
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.4830677290837 99.75 86.7330677290837 100 ;
		END PORT
	END pin_510
	PIN pin_511
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.16334661354585 99.75 86.41334661354585 100 ;
		END PORT
	END pin_511
	PIN pin_512
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.84362549800801 99.75 86.09362549800801 100 ;
		END PORT
	END pin_512
	PIN pin_513
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 85.52390438247016 99.75 85.77390438247016 100 ;
		END PORT
	END pin_513
	PIN pin_514
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.20418326693232 99.75 85.45418326693232 100 ;
		END PORT
	END pin_514
	PIN pin_515
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 84.88446215139447 99.75 85.13446215139447 100 ;
		END PORT
	END pin_515
	PIN pin_516
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 84.56474103585663 99.75 84.81474103585663 100 ;
		END PORT
	END pin_516
	PIN pin_517
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 84.24501992031878 99.75 84.49501992031878 100 ;
		END PORT
	END pin_517
	PIN pin_518
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.92529880478094 99.75 84.17529880478094 100 ;
		END PORT
	END pin_518
	PIN pin_519
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 83.60557768924309 99.75 83.85557768924309 100 ;
		END PORT
	END pin_519
	PIN pin_520
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 83.28585657370525 99.75 83.53585657370525 100 ;
		END PORT
	END pin_520
	PIN pin_521
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.9661354581674 99.75 83.2161354581674 100 ;
		END PORT
	END pin_521
	PIN pin_522
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.64641434262955 99.75 82.89641434262955 100 ;
		END PORT
	END pin_522
	PIN pin_523
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.32669322709171 99.75 82.57669322709171 100 ;
		END PORT
	END pin_523
	PIN pin_524
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.00697211155386 99.75 82.25697211155386 100 ;
		END PORT
	END pin_524
	PIN pin_525
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.68725099601602 99.75 81.93725099601602 100 ;
		END PORT
	END pin_525
	PIN pin_526
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 81.36752988047817 99.75 81.61752988047817 100 ;
		END PORT
	END pin_526
	PIN pin_527
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 81.04780876494033 99.75 81.29780876494033 100 ;
		END PORT
	END pin_527
	PIN pin_528
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 80.72808764940248 99.75 80.97808764940248 100 ;
		END PORT
	END pin_528
	PIN pin_529
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.40836653386464 99.75 80.65836653386464 100 ;
		END PORT
	END pin_529
	PIN pin_530
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.08864541832679 99.75 80.33864541832679 100 ;
		END PORT
	END pin_530
	PIN pin_531
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.76892430278895 99.75 80.01892430278895 100 ;
		END PORT
	END pin_531
	PIN pin_532
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.4492031872511 99.75 79.6992031872511 100 ;
		END PORT
	END pin_532
	PIN pin_533
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.12948207171326 99.75 79.37948207171326 100 ;
		END PORT
	END pin_533
	PIN pin_534
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 78.80976095617541 99.75 79.05976095617541 100 ;
		END PORT
	END pin_534
	PIN pin_535
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 78.49003984063756 99.75 78.74003984063756 100 ;
		END PORT
	END pin_535
	PIN pin_536
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 78.17031872509972 99.75 78.42031872509972 100 ;
		END PORT
	END pin_536
	PIN pin_537
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.85059760956187 99.75 78.10059760956187 100 ;
		END PORT
	END pin_537
	PIN pin_538
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 77.53087649402403 99.75 77.78087649402403 100 ;
		END PORT
	END pin_538
	PIN pin_539
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 77.21115537848618 99.75 77.46115537848618 100 ;
		END PORT
	END pin_539
	PIN pin_540
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 76.89143426294834 99.75 77.14143426294834 100 ;
		END PORT
	END pin_540
	PIN pin_541
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.57171314741049 99.75 76.82171314741049 100 ;
		END PORT
	END pin_541
	PIN pin_542
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.25199203187265 99.75 76.50199203187265 100 ;
		END PORT
	END pin_542
	PIN pin_543
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.9322709163348 99.75 76.1822709163348 100 ;
		END PORT
	END pin_543
	PIN pin_544
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 75.61254980079696 99.75 75.86254980079696 100 ;
		END PORT
	END pin_544
	PIN pin_545
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.29282868525911 99.75 75.54282868525911 100 ;
		END PORT
	END pin_545
	PIN pin_546
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.97310756972126 99.75 75.22310756972126 100 ;
		END PORT
	END pin_546
	PIN pin_547
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.65338645418342 99.75 74.90338645418342 100 ;
		END PORT
	END pin_547
	PIN pin_548
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 74.33366533864557 99.75 74.58366533864557 100 ;
		END PORT
	END pin_548
	PIN pin_549
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.01394422310773 99.75 74.26394422310773 100 ;
		END PORT
	END pin_549
	PIN pin_550
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 73.69422310756988 99.75 73.94422310756988 100 ;
		END PORT
	END pin_550
	PIN pin_551
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 73.37450199203204 99.75 73.62450199203204 100 ;
		END PORT
	END pin_551
	PIN pin_552
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 73.05478087649419 99.75 73.30478087649419 100 ;
		END PORT
	END pin_552
	PIN pin_553
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 72.73505976095635 99.75 72.98505976095635 100 ;
		END PORT
	END pin_553
	PIN pin_554
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 72.4153386454185 99.75 72.6653386454185 100 ;
		END PORT
	END pin_554
	PIN pin_555
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 72.09561752988066 99.75 72.34561752988066 100 ;
		END PORT
	END pin_555
	PIN pin_556
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 71.77589641434281 99.75 72.02589641434281 100 ;
		END PORT
	END pin_556
	PIN pin_557
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 71.45617529880496 99.75 71.70617529880496 100 ;
		END PORT
	END pin_557
	PIN pin_558
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 71.13645418326712 99.75 71.38645418326712 100 ;
		END PORT
	END pin_558
	PIN pin_559
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 70.81673306772927 99.75 71.06673306772927 100 ;
		END PORT
	END pin_559
	PIN pin_560
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.49701195219143 99.75 70.74701195219143 100 ;
		END PORT
	END pin_560
	PIN pin_561
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 70.17729083665358 99.75 70.42729083665358 100 ;
		END PORT
	END pin_561
	PIN pin_562
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 69.85756972111574 99.75 70.10756972111574 100 ;
		END PORT
	END pin_562
	PIN pin_563
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 69.53784860557789 99.75 69.78784860557789 100 ;
		END PORT
	END pin_563
	PIN pin_564
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 69.21812749004005 99.75 69.46812749004005 100 ;
		END PORT
	END pin_564
	PIN pin_565
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 68.8984063745022 99.75 69.1484063745022 100 ;
		END PORT
	END pin_565
	PIN pin_566
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 68.57868525896436 99.75 68.82868525896436 100 ;
		END PORT
	END pin_566
	PIN pin_567
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 68.25896414342651 99.75 68.50896414342651 100 ;
		END PORT
	END pin_567
	PIN pin_568
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 67.93924302788866 99.75 68.18924302788866 100 ;
		END PORT
	END pin_568
	PIN pin_569
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 67.61952191235082 99.75 67.86952191235082 100 ;
		END PORT
	END pin_569
	PIN pin_570
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.29980079681297 99.75 67.54980079681297 100 ;
		END PORT
	END pin_570
	PIN pin_571
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.98007968127513 99.75 67.23007968127513 100 ;
		END PORT
	END pin_571
	PIN pin_572
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.66035856573728 99.75 66.91035856573728 100 ;
		END PORT
	END pin_572
	PIN pin_573
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.34063745019944 99.75 66.59063745019944 100 ;
		END PORT
	END pin_573
	PIN pin_574
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.02091633466159 99.75 66.27091633466159 100 ;
		END PORT
	END pin_574
	PIN pin_575
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 65.70119521912375 99.75 65.95119521912375 100 ;
		END PORT
	END pin_575
	PIN pin_576
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 65.3814741035859 99.75 65.6314741035859 100 ;
		END PORT
	END pin_576
	PIN pin_577
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.06175298804806 99.75 65.31175298804806 100 ;
		END PORT
	END pin_577
	PIN pin_578
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 64.74203187251021 99.75 64.99203187251021 100 ;
		END PORT
	END pin_578
	PIN pin_579
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.42231075697237 99.75 64.67231075697237 100 ;
		END PORT
	END pin_579
	PIN pin_580
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 64.10258964143452 99.75 64.35258964143452 100 ;
		END PORT
	END pin_580
	PIN pin_581
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.782868525896674 99.75 64.03286852589667 100 ;
		END PORT
	END pin_581
	PIN pin_582
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.46314741035883 99.75 63.71314741035883 100 ;
		END PORT
	END pin_582
	PIN pin_583
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 63.14342629482098 99.75 63.39342629482098 100 ;
		END PORT
	END pin_583
	PIN pin_584
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.82370517928314 99.75 63.07370517928314 100 ;
		END PORT
	END pin_584
	PIN pin_585
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.50398406374529 99.75 62.75398406374529 100 ;
		END PORT
	END pin_585
	PIN pin_586
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 62.18426294820745 99.75 62.43426294820745 100 ;
		END PORT
	END pin_586
	PIN pin_587
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 61.8645418326696 99.75 62.1145418326696 100 ;
		END PORT
	END pin_587
	PIN pin_588
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 61.544820717131756 99.75 61.794820717131756 100 ;
		END PORT
	END pin_588
	PIN pin_589
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 61.22509960159391 99.75 61.47509960159391 100 ;
		END PORT
	END pin_589
	PIN pin_590
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 60.905378486056065 99.75 61.155378486056065 100 ;
		END PORT
	END pin_590
	PIN pin_591
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.58565737051822 99.75 60.83565737051822 100 ;
		END PORT
	END pin_591
	PIN pin_592
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.265936254980375 99.75 60.515936254980375 100 ;
		END PORT
	END pin_592
	PIN pin_593
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 59.94621513944253 99.75 60.19621513944253 100 ;
		END PORT
	END pin_593
	PIN pin_594
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 59.626494023904684 99.75 59.876494023904684 100 ;
		END PORT
	END pin_594
	PIN pin_595
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 59.30677290836684 99.75 59.55677290836684 100 ;
		END PORT
	END pin_595
	PIN pin_596
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.98705179282899 99.75 59.23705179282899 100 ;
		END PORT
	END pin_596
	PIN pin_597
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.66733067729115 99.75 58.91733067729115 100 ;
		END PORT
	END pin_597
	PIN pin_598
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.3476095617533 99.75 58.5976095617533 100 ;
		END PORT
	END pin_598
	PIN pin_599
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.02788844621546 99.75 58.27788844621546 100 ;
		END PORT
	END pin_599
	PIN pin_600
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.70816733067761 99.75 57.95816733067761 100 ;
		END PORT
	END pin_600
	PIN pin_601
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 57.388446215139766 99.75 57.638446215139766 100 ;
		END PORT
	END pin_601
	PIN pin_602
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.06872509960192 99.75 57.31872509960192 100 ;
		END PORT
	END pin_602
	PIN pin_603
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.749003984064075 99.75 56.999003984064075 100 ;
		END PORT
	END pin_603
	PIN pin_604
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 56.42928286852623 99.75 56.67928286852623 100 ;
		END PORT
	END pin_604
	PIN pin_605
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 56.109561752988384 99.75 56.359561752988384 100 ;
		END PORT
	END pin_605
	PIN pin_606
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.78984063745054 99.75 56.03984063745054 100 ;
		END PORT
	END pin_606
	PIN pin_607
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 55.47011952191269 99.75 55.72011952191269 100 ;
		END PORT
	END pin_607
	PIN pin_608
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.15039840637485 99.75 55.40039840637485 100 ;
		END PORT
	END pin_608
	PIN pin_609
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.830677290837 99.75 55.080677290837 100 ;
		END PORT
	END pin_609
	PIN pin_610
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 54.51095617529916 99.75 54.76095617529916 100 ;
		END PORT
	END pin_610
	PIN pin_611
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.19123505976131 99.75 54.44123505976131 100 ;
		END PORT
	END pin_611
	PIN pin_612
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.871513944223466 99.75 54.121513944223466 100 ;
		END PORT
	END pin_612
	PIN pin_613
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.55179282868562 99.75 53.80179282868562 100 ;
		END PORT
	END pin_613
	PIN pin_614
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 53.232071713147775 99.75 53.482071713147775 100 ;
		END PORT
	END pin_614
	PIN pin_615
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 52.91235059760993 99.75 53.16235059760993 100 ;
		END PORT
	END pin_615
	PIN pin_616
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 52.592629482072084 99.75 52.842629482072084 100 ;
		END PORT
	END pin_616
	PIN pin_617
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 52.27290836653424 99.75 52.52290836653424 100 ;
		END PORT
	END pin_617
	PIN pin_618
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 51.95318725099639 99.75 52.20318725099639 100 ;
		END PORT
	END pin_618
	PIN pin_619
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 51.63346613545855 99.75 51.88346613545855 100 ;
		END PORT
	END pin_619
	PIN pin_620
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.3137450199207 99.75 51.5637450199207 100 ;
		END PORT
	END pin_620
	PIN pin_621
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 50.99402390438286 99.75 51.24402390438286 100 ;
		END PORT
	END pin_621
	PIN pin_622
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.67430278884501 99.75 50.92430278884501 100 ;
		END PORT
	END pin_622
	PIN pin_623
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.354581673307166 99.75 50.604581673307166 100 ;
		END PORT
	END pin_623
	PIN pin_624
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.03486055776932 99.75 50.28486055776932 100 ;
		END PORT
	END pin_624
	PIN pin_625
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.715139442231475 99.75 49.965139442231475 100 ;
		END PORT
	END pin_625
	PIN pin_626
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.39541832669363 99.75 49.64541832669363 100 ;
		END PORT
	END pin_626
	PIN pin_627
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.075697211155784 99.75 49.325697211155784 100 ;
		END PORT
	END pin_627
	PIN pin_628
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.75597609561794 99.75 49.00597609561794 100 ;
		END PORT
	END pin_628
	PIN pin_629
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.43625498008009 99.75 48.68625498008009 100 ;
		END PORT
	END pin_629
	PIN pin_630
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 48.11653386454225 99.75 48.36653386454225 100 ;
		END PORT
	END pin_630
	PIN pin_631
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 47.7968127490044 99.75 48.0468127490044 100 ;
		END PORT
	END pin_631
	PIN pin_632
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.47709163346656 99.75 47.72709163346656 100 ;
		END PORT
	END pin_632
	PIN pin_633
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 47.15737051792871 99.75 47.40737051792871 100 ;
		END PORT
	END pin_633
	PIN pin_634
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.837649402390866 99.75 47.087649402390866 100 ;
		END PORT
	END pin_634
	PIN pin_635
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 46.51792828685302 99.75 46.76792828685302 100 ;
		END PORT
	END pin_635
	PIN pin_636
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 46.198207171315175 99.75 46.448207171315175 100 ;
		END PORT
	END pin_636
	PIN pin_637
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.87848605577733 99.75 46.12848605577733 100 ;
		END PORT
	END pin_637
	PIN pin_638
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 45.558764940239485 99.75 45.808764940239485 100 ;
		END PORT
	END pin_638
	PIN pin_639
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.23904382470164 99.75 45.48904382470164 100 ;
		END PORT
	END pin_639
	PIN pin_640
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.919322709163794 99.75 45.169322709163794 100 ;
		END PORT
	END pin_640
	PIN pin_641
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.59960159362595 99.75 44.84960159362595 100 ;
		END PORT
	END pin_641
	PIN pin_642
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 44.2798804780881 99.75 44.5298804780881 100 ;
		END PORT
	END pin_642
	PIN pin_643
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 43.96015936255026 99.75 44.21015936255026 100 ;
		END PORT
	END pin_643
	PIN pin_644
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.64043824701241 99.75 43.89043824701241 100 ;
		END PORT
	END pin_644
	PIN pin_645
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 43.32071713147457 99.75 43.57071713147457 100 ;
		END PORT
	END pin_645
	PIN pin_646
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 43.00099601593672 99.75 43.25099601593672 100 ;
		END PORT
	END pin_646
	PIN pin_647
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.681274900398876 99.75 42.931274900398876 100 ;
		END PORT
	END pin_647
	PIN pin_648
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 42.36155378486103 99.75 42.61155378486103 100 ;
		END PORT
	END pin_648
	PIN pin_649
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 42.041832669323185 99.75 42.291832669323185 100 ;
		END PORT
	END pin_649
	PIN pin_650
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 41.72211155378534 99.75 41.97211155378534 100 ;
		END PORT
	END pin_650
	PIN pin_651
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.402390438247494 99.75 41.652390438247494 100 ;
		END PORT
	END pin_651
	PIN pin_652
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.08266932270965 99.75 41.33266932270965 100 ;
		END PORT
	END pin_652
	PIN pin_653
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.7629482071718 99.75 41.0129482071718 100 ;
		END PORT
	END pin_653
	PIN pin_654
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.44322709163396 99.75 40.69322709163396 100 ;
		END PORT
	END pin_654
	PIN pin_655
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 40.12350597609611 99.75 40.37350597609611 100 ;
		END PORT
	END pin_655
	PIN pin_656
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 39.80378486055827 99.75 40.05378486055827 100 ;
		END PORT
	END pin_656
	PIN pin_657
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 39.48406374502042 99.75 39.73406374502042 100 ;
		END PORT
	END pin_657
	PIN pin_658
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 39.164342629482576 99.75 39.414342629482576 100 ;
		END PORT
	END pin_658
	PIN pin_659
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 38.84462151394473 99.75 39.09462151394473 100 ;
		END PORT
	END pin_659
	PIN pin_660
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.524900398406885 99.75 38.774900398406885 100 ;
		END PORT
	END pin_660
	PIN pin_661
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 38.20517928286904 99.75 38.45517928286904 100 ;
		END PORT
	END pin_661
	PIN pin_662
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 37.885458167331194 99.75 38.135458167331194 100 ;
		END PORT
	END pin_662
	PIN pin_663
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 37.56573705179335 99.75 37.81573705179335 100 ;
		END PORT
	END pin_663
	PIN pin_664
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.2460159362555 99.75 37.4960159362555 100 ;
		END PORT
	END pin_664
	PIN pin_665
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 36.92629482071766 99.75 37.17629482071766 100 ;
		END PORT
	END pin_665
	PIN pin_666
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.60657370517981 99.75 36.85657370517981 100 ;
		END PORT
	END pin_666
	PIN pin_667
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.28685258964197 99.75 36.53685258964197 100 ;
		END PORT
	END pin_667
	PIN pin_668
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.96713147410412 99.75 36.21713147410412 100 ;
		END PORT
	END pin_668
	PIN pin_669
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 35.647410358566276 99.75 35.897410358566276 100 ;
		END PORT
	END pin_669
	PIN pin_670
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 35.32768924302843 99.75 35.57768924302843 100 ;
		END PORT
	END pin_670
	PIN pin_671
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 35.007968127490585 99.75 35.257968127490585 100 ;
		END PORT
	END pin_671
	PIN pin_672
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.68824701195274 99.75 34.93824701195274 100 ;
		END PORT
	END pin_672
	PIN pin_673
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.368525896414894 99.75 34.618525896414894 100 ;
		END PORT
	END pin_673
	PIN pin_674
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 34.04880478087705 99.75 34.29880478087705 100 ;
		END PORT
	END pin_674
	PIN pin_675
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.7290836653392 99.75 33.9790836653392 100 ;
		END PORT
	END pin_675
	PIN pin_676
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.40936254980136 99.75 33.65936254980136 100 ;
		END PORT
	END pin_676
	PIN pin_677
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 33.08964143426351 99.75 33.33964143426351 100 ;
		END PORT
	END pin_677
	PIN pin_678
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 32.76992031872567 99.75 33.01992031872567 100 ;
		END PORT
	END pin_678
	PIN pin_679
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 32.45019920318782 99.75 32.70019920318782 100 ;
		END PORT
	END pin_679
	PIN pin_680
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.130478087649976 99.75 32.380478087649976 100 ;
		END PORT
	END pin_680
	PIN pin_681
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.81075697211213 99.75 32.06075697211213 100 ;
		END PORT
	END pin_681
	PIN pin_682
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 31.491035856574282 99.75 31.741035856574282 100 ;
		END PORT
	END pin_682
	PIN pin_683
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 31.171314741036433 99.75 31.421314741036433 100 ;
		END PORT
	END pin_683
	PIN pin_684
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.851593625498584 99.75 31.101593625498584 100 ;
		END PORT
	END pin_684
	PIN pin_685
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 30.531872509960735 99.75 30.781872509960735 100 ;
		END PORT
	END pin_685
	PIN pin_686
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 30.212151394422886 99.75 30.462151394422886 100 ;
		END PORT
	END pin_686
	PIN pin_687
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.892430278885037 99.75 30.142430278885037 100 ;
		END PORT
	END pin_687
	PIN pin_688
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 29.572709163347188 99.75 29.822709163347188 100 ;
		END PORT
	END pin_688
	PIN pin_689
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 29.25298804780934 99.75 29.50298804780934 100 ;
		END PORT
	END pin_689
	PIN pin_690
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 28.93326693227149 99.75 29.18326693227149 100 ;
		END PORT
	END pin_690
	PIN pin_691
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.61354581673364 99.75 28.86354581673364 100 ;
		END PORT
	END pin_691
	PIN pin_692
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 28.293824701195792 99.75 28.543824701195792 100 ;
		END PORT
	END pin_692
	PIN pin_693
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.974103585657943 99.75 28.224103585657943 100 ;
		END PORT
	END pin_693
	PIN pin_694
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.654382470120094 99.75 27.904382470120094 100 ;
		END PORT
	END pin_694
	PIN pin_695
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.334661354582245 99.75 27.584661354582245 100 ;
		END PORT
	END pin_695
	PIN pin_696
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.014940239044396 99.75 27.264940239044396 100 ;
		END PORT
	END pin_696
	PIN pin_697
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.695219123506547 99.75 26.945219123506547 100 ;
		END PORT
	END pin_697
	PIN pin_698
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 26.375498007968698 99.75 26.625498007968698 100 ;
		END PORT
	END pin_698
	PIN pin_699
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.05577689243085 99.75 26.30577689243085 100 ;
		END PORT
	END pin_699
	PIN pin_700
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 25.736055776893 99.75 25.986055776893 100 ;
		END PORT
	END pin_700
	PIN pin_701
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 25.41633466135515 99.75 25.66633466135515 100 ;
		END PORT
	END pin_701
	PIN pin_702
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 25.096613545817302 99.75 25.346613545817302 100 ;
		END PORT
	END pin_702
	PIN pin_703
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 24.776892430279453 99.75 25.026892430279453 100 ;
		END PORT
	END pin_703
	PIN pin_704
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.457171314741604 99.75 24.707171314741604 100 ;
		END PORT
	END pin_704
	PIN pin_705
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 24.137450199203755 99.75 24.387450199203755 100 ;
		END PORT
	END pin_705
	PIN pin_706
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.817729083665906 99.75 24.067729083665906 100 ;
		END PORT
	END pin_706
	PIN pin_707
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 23.498007968128057 99.75 23.748007968128057 100 ;
		END PORT
	END pin_707
	PIN pin_708
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 23.178286852590208 99.75 23.428286852590208 100 ;
		END PORT
	END pin_708
	PIN pin_709
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.85856573705236 99.75 23.10856573705236 100 ;
		END PORT
	END pin_709
	PIN pin_710
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 22.53884462151451 99.75 22.78884462151451 100 ;
		END PORT
	END pin_710
	PIN pin_711
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.21912350597666 99.75 22.46912350597666 100 ;
		END PORT
	END pin_711
	PIN pin_712
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.899402390438812 99.75 22.149402390438812 100 ;
		END PORT
	END pin_712
	PIN pin_713
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 21.579681274900963 99.75 21.829681274900963 100 ;
		END PORT
	END pin_713
	PIN pin_714
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.259960159363114 99.75 21.509960159363114 100 ;
		END PORT
	END pin_714
	PIN pin_715
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 20.940239043825265 99.75 21.190239043825265 100 ;
		END PORT
	END pin_715
	PIN pin_716
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 20.620517928287416 99.75 20.870517928287416 100 ;
		END PORT
	END pin_716
	PIN pin_717
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 20.300796812749567 99.75 20.550796812749567 100 ;
		END PORT
	END pin_717
	PIN pin_718
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.98107569721172 99.75 20.23107569721172 100 ;
		END PORT
	END pin_718
	PIN pin_719
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 19.66135458167387 99.75 19.91135458167387 100 ;
		END PORT
	END pin_719
	PIN pin_720
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.34163346613602 99.75 19.59163346613602 100 ;
		END PORT
	END pin_720
	PIN pin_721
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.02191235059817 99.75 19.27191235059817 100 ;
		END PORT
	END pin_721
	PIN pin_722
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 18.702191235060322 99.75 18.952191235060322 100 ;
		END PORT
	END pin_722
	PIN pin_723
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 18.382470119522473 99.75 18.632470119522473 100 ;
		END PORT
	END pin_723
	PIN pin_724
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.062749003984624 99.75 18.312749003984624 100 ;
		END PORT
	END pin_724
	PIN pin_725
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 17.743027888446775 99.75 17.993027888446775 100 ;
		END PORT
	END pin_725
	PIN pin_726
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 17.423306772908926 99.75 17.673306772908926 100 ;
		END PORT
	END pin_726
	PIN pin_727
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.103585657371077 99.75 17.353585657371077 100 ;
		END PORT
	END pin_727
	PIN pin_728
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.78386454183323 99.75 17.03386454183323 100 ;
		END PORT
	END pin_728
	PIN pin_729
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.46414342629538 99.75 16.71414342629538 100 ;
		END PORT
	END pin_729
	PIN pin_730
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.14442231075753 99.75 16.39442231075753 100 ;
		END PORT
	END pin_730
	PIN pin_731
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.824701195219681 99.75 16.07470119521968 100 ;
		END PORT
	END pin_731
	PIN pin_732
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 15.504980079681832 99.75 15.754980079681832 100 ;
		END PORT
	END pin_732
	PIN pin_733
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 15.185258964143983 99.75 15.435258964143983 100 ;
		END PORT
	END pin_733
	PIN pin_734
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.865537848606134 99.75 15.115537848606134 100 ;
		END PORT
	END pin_734
	PIN pin_735
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 14.545816733068285 99.75 14.795816733068285 100 ;
		END PORT
	END pin_735
	PIN pin_736
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.226095617530436 99.75 14.476095617530436 100 ;
		END PORT
	END pin_736
	PIN pin_737
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 13.906374501992588 99.75 14.156374501992588 100 ;
		END PORT
	END pin_737
	PIN pin_738
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 13.586653386454739 99.75 13.836653386454739 100 ;
		END PORT
	END pin_738
	PIN pin_739
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 13.26693227091689 99.75 13.51693227091689 100 ;
		END PORT
	END pin_739
	PIN pin_740
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 12.94721115537904 99.75 13.19721115537904 100 ;
		END PORT
	END pin_740
	PIN pin_741
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 12.627490039841192 99.75 12.877490039841192 100 ;
		END PORT
	END pin_741
	PIN pin_742
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 12.307768924303343 99.75 12.557768924303343 100 ;
		END PORT
	END pin_742
	PIN pin_743
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 11.988047808765494 99.75 12.238047808765494 100 ;
		END PORT
	END pin_743
	PIN pin_744
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 11.668326693227645 99.75 11.918326693227645 100 ;
		END PORT
	END pin_744
	PIN pin_745
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.348605577689796 99.75 11.598605577689796 100 ;
		END PORT
	END pin_745
	PIN pin_746
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.028884462151947 99.75 11.278884462151947 100 ;
		END PORT
	END pin_746
	PIN pin_747
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 10.709163346614098 99.75 10.959163346614098 100 ;
		END PORT
	END pin_747
	PIN pin_748
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 10.389442231076249 99.75 10.639442231076249 100 ;
		END PORT
	END pin_748
	PIN pin_749
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 10.0697211155384 99.75 10.3197211155384 100 ;
		END PORT
	END pin_749
	PIN pin_750
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 10.069721115537849 0 10.319721115537849 0.25 ;
		END PORT
	END pin_750
	PIN pin_751
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 10.389442231075698 0 10.639442231075698 0.25 ;
		END PORT
	END pin_751
	PIN pin_752
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 10.709163346613547 0 10.959163346613547 0.25 ;
		END PORT
	END pin_752
	PIN pin_753
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.028884462151396 0 11.278884462151396 0.25 ;
		END PORT
	END pin_753
	PIN pin_754
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.348605577689245 0 11.598605577689245 0.25 ;
		END PORT
	END pin_754
	PIN pin_755
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.668326693227094 0 11.918326693227094 0.25 ;
		END PORT
	END pin_755
	PIN pin_756
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 11.988047808764943 0 12.238047808764943 0.25 ;
		END PORT
	END pin_756
	PIN pin_757
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 12.307768924302792 0 12.557768924302792 0.25 ;
		END PORT
	END pin_757
	PIN pin_758
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 12.627490039840641 0 12.877490039840641 0.25 ;
		END PORT
	END pin_758
	PIN pin_759
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 12.94721115537849 0 13.19721115537849 0.25 ;
		END PORT
	END pin_759
	PIN pin_760
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 13.266932270916339 0 13.516932270916339 0.25 ;
		END PORT
	END pin_760
	PIN pin_761
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 13.586653386454188 0 13.836653386454188 0.25 ;
		END PORT
	END pin_761
	PIN pin_762
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 13.906374501992037 0 14.156374501992037 0.25 ;
		END PORT
	END pin_762
	PIN pin_763
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 14.226095617529886 0 14.476095617529886 0.25 ;
		END PORT
	END pin_763
	PIN pin_764
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.545816733067735 0 14.795816733067735 0.25 ;
		END PORT
	END pin_764
	PIN pin_765
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 14.865537848605584 0 15.115537848605584 0.25 ;
		END PORT
	END pin_765
	PIN pin_766
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 15.185258964143433 0 15.435258964143433 0.25 ;
		END PORT
	END pin_766
	PIN pin_767
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.504980079681282 0 15.754980079681282 0.25 ;
		END PORT
	END pin_767
	PIN pin_768
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 15.82470119521913 0 16.07470119521913 0.25 ;
		END PORT
	END pin_768
	PIN pin_769
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 16.14442231075698 0 16.39442231075698 0.25 ;
		END PORT
	END pin_769
	PIN pin_770
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 16.46414342629483 0 16.71414342629483 0.25 ;
		END PORT
	END pin_770
	PIN pin_771
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 16.783864541832678 0 17.033864541832678 0.25 ;
		END PORT
	END pin_771
	PIN pin_772
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 17.103585657370527 0 17.353585657370527 0.25 ;
		END PORT
	END pin_772
	PIN pin_773
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 17.423306772908376 0 17.673306772908376 0.25 ;
		END PORT
	END pin_773
	PIN pin_774
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 17.743027888446225 0 17.993027888446225 0.25 ;
		END PORT
	END pin_774
	PIN pin_775
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.062749003984074 0 18.312749003984074 0.25 ;
		END PORT
	END pin_775
	PIN pin_776
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 18.382470119521923 0 18.632470119521923 0.25 ;
		END PORT
	END pin_776
	PIN pin_777
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.70219123505977 0 18.95219123505977 0.25 ;
		END PORT
	END pin_777
	PIN pin_778
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.02191235059762 0 19.27191235059762 0.25 ;
		END PORT
	END pin_778
	PIN pin_779
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.34163346613547 0 19.59163346613547 0.25 ;
		END PORT
	END pin_779
	PIN pin_780
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.66135458167332 0 19.91135458167332 0.25 ;
		END PORT
	END pin_780
	PIN pin_781
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 19.981075697211168 0 20.231075697211168 0.25 ;
		END PORT
	END pin_781
	PIN pin_782
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.300796812749017 0 20.550796812749017 0.25 ;
		END PORT
	END pin_782
	PIN pin_783
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 20.620517928286866 0 20.870517928286866 0.25 ;
		END PORT
	END pin_783
	PIN pin_784
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 20.940239043824715 0 21.190239043824715 0.25 ;
		END PORT
	END pin_784
	PIN pin_785
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 21.259960159362564 0 21.509960159362564 0.25 ;
		END PORT
	END pin_785
	PIN pin_786
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.579681274900413 0 21.829681274900413 0.25 ;
		END PORT
	END pin_786
	PIN pin_787
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 21.89940239043826 0 22.14940239043826 0.25 ;
		END PORT
	END pin_787
	PIN pin_788
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 22.21912350597611 0 22.46912350597611 0.25 ;
		END PORT
	END pin_788
	PIN pin_789
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 22.53884462151396 0 22.78884462151396 0.25 ;
		END PORT
	END pin_789
	PIN pin_790
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 22.85856573705181 0 23.10856573705181 0.25 ;
		END PORT
	END pin_790
	PIN pin_791
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 23.178286852589657 0 23.428286852589657 0.25 ;
		END PORT
	END pin_791
	PIN pin_792
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 23.498007968127506 0 23.748007968127506 0.25 ;
		END PORT
	END pin_792
	PIN pin_793
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 23.817729083665355 0 24.067729083665355 0.25 ;
		END PORT
	END pin_793
	PIN pin_794
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.137450199203204 0 24.387450199203204 0.25 ;
		END PORT
	END pin_794
	PIN pin_795
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 24.457171314741053 0 24.707171314741053 0.25 ;
		END PORT
	END pin_795
	PIN pin_796
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 24.776892430278902 0 25.026892430278902 0.25 ;
		END PORT
	END pin_796
	PIN pin_797
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 25.09661354581675 0 25.34661354581675 0.25 ;
		END PORT
	END pin_797
	PIN pin_798
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 25.4163346613546 0 25.6663346613546 0.25 ;
		END PORT
	END pin_798
	PIN pin_799
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 25.73605577689245 0 25.98605577689245 0.25 ;
		END PORT
	END pin_799
	PIN pin_800
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.0557768924303 0 26.3057768924303 0.25 ;
		END PORT
	END pin_800
	PIN pin_801
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 26.375498007968147 0 26.625498007968147 0.25 ;
		END PORT
	END pin_801
	PIN pin_802
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 26.695219123505996 0 26.945219123505996 0.25 ;
		END PORT
	END pin_802
	PIN pin_803
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 27.014940239043845 0 27.264940239043845 0.25 ;
		END PORT
	END pin_803
	PIN pin_804
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 27.334661354581694 0 27.584661354581694 0.25 ;
		END PORT
	END pin_804
	PIN pin_805
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 27.654382470119543 0 27.904382470119543 0.25 ;
		END PORT
	END pin_805
	PIN pin_806
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 27.974103585657392 0 28.224103585657392 0.25 ;
		END PORT
	END pin_806
	PIN pin_807
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.29382470119524 0 28.54382470119524 0.25 ;
		END PORT
	END pin_807
	PIN pin_808
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 28.61354581673309 0 28.86354581673309 0.25 ;
		END PORT
	END pin_808
	PIN pin_809
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 28.93326693227094 0 29.18326693227094 0.25 ;
		END PORT
	END pin_809
	PIN pin_810
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 29.25298804780879 0 29.50298804780879 0.25 ;
		END PORT
	END pin_810
	PIN pin_811
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 29.572709163346637 0 29.822709163346637 0.25 ;
		END PORT
	END pin_811
	PIN pin_812
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 29.892430278884486 0 30.142430278884486 0.25 ;
		END PORT
	END pin_812
	PIN pin_813
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 30.212151394422335 0 30.462151394422335 0.25 ;
		END PORT
	END pin_813
	PIN pin_814
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 30.531872509960184 0 30.781872509960184 0.25 ;
		END PORT
	END pin_814
	PIN pin_815
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 30.851593625498033 0 31.101593625498033 0.25 ;
		END PORT
	END pin_815
	PIN pin_816
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.171314741035882 0 31.421314741035882 0.25 ;
		END PORT
	END pin_816
	PIN pin_817
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 31.49103585657373 0 31.74103585657373 0.25 ;
		END PORT
	END pin_817
	PIN pin_818
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 31.81075697211158 0 32.06075697211158 0.25 ;
		END PORT
	END pin_818
	PIN pin_819
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 32.13047808764942 0 32.38047808764942 0.25 ;
		END PORT
	END pin_819
	PIN pin_820
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.45019920318727 0 32.70019920318727 0.25 ;
		END PORT
	END pin_820
	PIN pin_821
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.76992031872511 0 33.01992031872511 0.25 ;
		END PORT
	END pin_821
	PIN pin_822
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.08964143426296 0 33.33964143426296 0.25 ;
		END PORT
	END pin_822
	PIN pin_823
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.409362549800804 0 33.659362549800804 0.25 ;
		END PORT
	END pin_823
	PIN pin_824
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 33.72908366533865 0 33.97908366533865 0.25 ;
		END PORT
	END pin_824
	PIN pin_825
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 34.048804780876495 0 34.298804780876495 0.25 ;
		END PORT
	END pin_825
	PIN pin_826
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 34.36852589641434 0 34.61852589641434 0.25 ;
		END PORT
	END pin_826
	PIN pin_827
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 34.688247011952186 0 34.938247011952186 0.25 ;
		END PORT
	END pin_827
	PIN pin_828
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.00796812749003 0 35.25796812749003 0.25 ;
		END PORT
	END pin_828
	PIN pin_829
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 35.327689243027876 0 35.577689243027876 0.25 ;
		END PORT
	END pin_829
	PIN pin_830
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 35.64741035856572 0 35.89741035856572 0.25 ;
		END PORT
	END pin_830
	PIN pin_831
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.96713147410357 0 36.21713147410357 0.25 ;
		END PORT
	END pin_831
	PIN pin_832
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.28685258964141 0 36.53685258964141 0.25 ;
		END PORT
	END pin_832
	PIN pin_833
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.60657370517926 0 36.85657370517926 0.25 ;
		END PORT
	END pin_833
	PIN pin_834
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 36.926294820717104 0 37.176294820717104 0.25 ;
		END PORT
	END pin_834
	PIN pin_835
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.24601593625495 0 37.49601593625495 0.25 ;
		END PORT
	END pin_835
	PIN pin_836
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 37.565737051792794 0 37.815737051792794 0.25 ;
		END PORT
	END pin_836
	PIN pin_837
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 37.88545816733064 0 38.13545816733064 0.25 ;
		END PORT
	END pin_837
	PIN pin_838
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 38.205179282868485 0 38.455179282868485 0.25 ;
		END PORT
	END pin_838
	PIN pin_839
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 38.52490039840633 0 38.77490039840633 0.25 ;
		END PORT
	END pin_839
	PIN pin_840
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 38.844621513944176 0 39.094621513944176 0.25 ;
		END PORT
	END pin_840
	PIN pin_841
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 39.16434262948202 0 39.41434262948202 0.25 ;
		END PORT
	END pin_841
	PIN pin_842
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 39.48406374501987 0 39.73406374501987 0.25 ;
		END PORT
	END pin_842
	PIN pin_843
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 39.80378486055771 0 40.05378486055771 0.25 ;
		END PORT
	END pin_843
	PIN pin_844
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 40.12350597609556 0 40.37350597609556 0.25 ;
		END PORT
	END pin_844
	PIN pin_845
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 40.4432270916334 0 40.6932270916334 0.25 ;
		END PORT
	END pin_845
	PIN pin_846
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.76294820717125 0 41.01294820717125 0.25 ;
		END PORT
	END pin_846
	PIN pin_847
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.082669322709094 0 41.332669322709094 0.25 ;
		END PORT
	END pin_847
	PIN pin_848
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 41.40239043824694 0 41.65239043824694 0.25 ;
		END PORT
	END pin_848
	PIN pin_849
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 41.722111553784785 0 41.972111553784785 0.25 ;
		END PORT
	END pin_849
	PIN pin_850
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 42.04183266932263 0 42.29183266932263 0.25 ;
		END PORT
	END pin_850
	PIN pin_851
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 42.361553784860476 0 42.611553784860476 0.25 ;
		END PORT
	END pin_851
	PIN pin_852
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 42.68127490039832 0 42.93127490039832 0.25 ;
		END PORT
	END pin_852
	PIN pin_853
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 43.00099601593617 0 43.25099601593617 0.25 ;
		END PORT
	END pin_853
	PIN pin_854
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 43.32071713147401 0 43.57071713147401 0.25 ;
		END PORT
	END pin_854
	PIN pin_855
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 43.64043824701186 0 43.89043824701186 0.25 ;
		END PORT
	END pin_855
	PIN pin_856
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 43.9601593625497 0 44.2101593625497 0.25 ;
		END PORT
	END pin_856
	PIN pin_857
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.27988047808755 0 44.52988047808755 0.25 ;
		END PORT
	END pin_857
	PIN pin_858
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 44.599601593625394 0 44.849601593625394 0.25 ;
		END PORT
	END pin_858
	PIN pin_859
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.91932270916324 0 45.16932270916324 0.25 ;
		END PORT
	END pin_859
	PIN pin_860
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 45.239043824701085 0 45.489043824701085 0.25 ;
		END PORT
	END pin_860
	PIN pin_861
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 45.55876494023893 0 45.80876494023893 0.25 ;
		END PORT
	END pin_861
	PIN pin_862
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 45.878486055776776 0 46.128486055776776 0.25 ;
		END PORT
	END pin_862
	PIN pin_863
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 46.19820717131462 0 46.44820717131462 0.25 ;
		END PORT
	END pin_863
	PIN pin_864
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 46.51792828685247 0 46.76792828685247 0.25 ;
		END PORT
	END pin_864
	PIN pin_865
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 46.83764940239031 0 47.08764940239031 0.25 ;
		END PORT
	END pin_865
	PIN pin_866
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.15737051792816 0 47.40737051792816 0.25 ;
		END PORT
	END pin_866
	PIN pin_867
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.477091633466 0 47.727091633466 0.25 ;
		END PORT
	END pin_867
	PIN pin_868
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 47.79681274900385 0 48.04681274900385 0.25 ;
		END PORT
	END pin_868
	PIN pin_869
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 48.116533864541694 0 48.366533864541694 0.25 ;
		END PORT
	END pin_869
	PIN pin_870
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 48.43625498007954 0 48.68625498007954 0.25 ;
		END PORT
	END pin_870
	PIN pin_871
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 48.755976095617385 0 49.005976095617385 0.25 ;
		END PORT
	END pin_871
	PIN pin_872
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.07569721115523 0 49.32569721115523 0.25 ;
		END PORT
	END pin_872
	PIN pin_873
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 49.395418326693076 0 49.645418326693076 0.25 ;
		END PORT
	END pin_873
	PIN pin_874
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.71513944223092 0 49.96513944223092 0.25 ;
		END PORT
	END pin_874
	PIN pin_875
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.034860557768766 0 50.284860557768766 0.25 ;
		END PORT
	END pin_875
	PIN pin_876
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 50.35458167330661 0 50.60458167330661 0.25 ;
		END PORT
	END pin_876
	PIN pin_877
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 50.67430278884446 0 50.92430278884446 0.25 ;
		END PORT
	END pin_877
	PIN pin_878
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.9940239043823 0 51.2440239043823 0.25 ;
		END PORT
	END pin_878
	PIN pin_879
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 51.31374501992015 0 51.56374501992015 0.25 ;
		END PORT
	END pin_879
	PIN pin_880
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 51.633466135457994 0 51.883466135457994 0.25 ;
		END PORT
	END pin_880
	PIN pin_881
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 51.95318725099584 0 52.20318725099584 0.25 ;
		END PORT
	END pin_881
	PIN pin_882
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 52.272908366533684 0 52.522908366533684 0.25 ;
		END PORT
	END pin_882
	PIN pin_883
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 52.59262948207153 0 52.84262948207153 0.25 ;
		END PORT
	END pin_883
	PIN pin_884
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 52.912350597609375 0 53.162350597609375 0.25 ;
		END PORT
	END pin_884
	PIN pin_885
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 53.23207171314722 0 53.48207171314722 0.25 ;
		END PORT
	END pin_885
	PIN pin_886
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 53.551792828685066 0 53.801792828685066 0.25 ;
		END PORT
	END pin_886
	PIN pin_887
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 53.87151394422291 0 54.12151394422291 0.25 ;
		END PORT
	END pin_887
	PIN pin_888
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 54.19123505976076 0 54.44123505976076 0.25 ;
		END PORT
	END pin_888
	PIN pin_889
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.5109561752986 0 54.7609561752986 0.25 ;
		END PORT
	END pin_889
	PIN pin_890
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 54.83067729083645 0 55.08067729083645 0.25 ;
		END PORT
	END pin_890
	PIN pin_891
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.15039840637429 0 55.40039840637429 0.25 ;
		END PORT
	END pin_891
	PIN pin_892
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.47011952191214 0 55.72011952191214 0.25 ;
		END PORT
	END pin_892
	PIN pin_893
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.789840637449984 0 56.039840637449984 0.25 ;
		END PORT
	END pin_893
	PIN pin_894
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 56.10956175298783 0 56.35956175298783 0.25 ;
		END PORT
	END pin_894
	PIN pin_895
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.429282868525675 0 56.679282868525675 0.25 ;
		END PORT
	END pin_895
	PIN pin_896
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 56.74900398406352 0 56.99900398406352 0.25 ;
		END PORT
	END pin_896
	PIN pin_897
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.068725099601366 0 57.318725099601366 0.25 ;
		END PORT
	END pin_897
	PIN pin_898
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 57.38844621513921 0 57.63844621513921 0.25 ;
		END PORT
	END pin_898
	PIN pin_899
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.70816733067706 0 57.95816733067706 0.25 ;
		END PORT
	END pin_899
	PIN pin_900
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.0278884462149 0 58.2778884462149 0.25 ;
		END PORT
	END pin_900
	PIN pin_901
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 58.34760956175275 0 58.59760956175275 0.25 ;
		END PORT
	END pin_901
	PIN pin_902
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 58.66733067729059 0 58.91733067729059 0.25 ;
		END PORT
	END pin_902
	PIN pin_903
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.98705179282844 0 59.23705179282844 0.25 ;
		END PORT
	END pin_903
	PIN pin_904
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 59.306772908366284 0 59.556772908366284 0.25 ;
		END PORT
	END pin_904
	PIN pin_905
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 59.62649402390413 0 59.87649402390413 0.25 ;
		END PORT
	END pin_905
	PIN pin_906
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 59.946215139441975 0 60.196215139441975 0.25 ;
		END PORT
	END pin_906
	PIN pin_907
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 60.26593625497982 0 60.51593625497982 0.25 ;
		END PORT
	END pin_907
	PIN pin_908
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 60.585657370517666 0 60.835657370517666 0.25 ;
		END PORT
	END pin_908
	PIN pin_909
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 60.90537848605551 0 61.15537848605551 0.25 ;
		END PORT
	END pin_909
	PIN pin_910
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 61.22509960159336 0 61.47509960159336 0.25 ;
		END PORT
	END pin_910
	PIN pin_911
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 61.5448207171312 0 61.7948207171312 0.25 ;
		END PORT
	END pin_911
	PIN pin_912
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 61.86454183266905 0 62.11454183266905 0.25 ;
		END PORT
	END pin_912
	PIN pin_913
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 62.18426294820689 0 62.43426294820689 0.25 ;
		END PORT
	END pin_913
	PIN pin_914
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.50398406374474 0 62.75398406374474 0.25 ;
		END PORT
	END pin_914
	PIN pin_915
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.823705179282584 0 63.073705179282584 0.25 ;
		END PORT
	END pin_915
	PIN pin_916
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.14342629482043 0 63.39342629482043 0.25 ;
		END PORT
	END pin_916
	PIN pin_917
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.463147410358275 0 63.713147410358275 0.25 ;
		END PORT
	END pin_917
	PIN pin_918
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.78286852589612 0 64.03286852589612 0.25 ;
		END PORT
	END pin_918
	PIN pin_919
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 64.10258964143397 0 64.35258964143397 0.25 ;
		END PORT
	END pin_919
	PIN pin_920
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 64.42231075697181 0 64.67231075697181 0.25 ;
		END PORT
	END pin_920
	PIN pin_921
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 64.74203187250966 0 64.99203187250966 0.25 ;
		END PORT
	END pin_921
	PIN pin_922
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.0617529880475 0 65.3117529880475 0.25 ;
		END PORT
	END pin_922
	PIN pin_923
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.38147410358535 0 65.63147410358535 0.25 ;
		END PORT
	END pin_923
	PIN pin_924
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 65.70119521912319 0 65.95119521912319 0.25 ;
		END PORT
	END pin_924
	PIN pin_925
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.02091633466104 0 66.27091633466104 0.25 ;
		END PORT
	END pin_925
	PIN pin_926
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.34063745019888 0 66.59063745019888 0.25 ;
		END PORT
	END pin_926
	PIN pin_927
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 66.66035856573673 0 66.91035856573673 0.25 ;
		END PORT
	END pin_927
	PIN pin_928
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 66.98007968127457 0 67.23007968127457 0.25 ;
		END PORT
	END pin_928
	PIN pin_929
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.29980079681242 0 67.54980079681242 0.25 ;
		END PORT
	END pin_929
	PIN pin_930
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 67.61952191235027 0 67.86952191235027 0.25 ;
		END PORT
	END pin_930
	PIN pin_931
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 67.93924302788811 0 68.18924302788811 0.25 ;
		END PORT
	END pin_931
	PIN pin_932
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 68.25896414342596 0 68.50896414342596 0.25 ;
		END PORT
	END pin_932
	PIN pin_933
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 68.5786852589638 0 68.8286852589638 0.25 ;
		END PORT
	END pin_933
	PIN pin_934
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 68.89840637450165 0 69.14840637450165 0.25 ;
		END PORT
	END pin_934
	PIN pin_935
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 69.21812749003949 0 69.46812749003949 0.25 ;
		END PORT
	END pin_935
	PIN pin_936
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 69.53784860557734 0 69.78784860557734 0.25 ;
		END PORT
	END pin_936
	PIN pin_937
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 69.85756972111518 0 70.10756972111518 0.25 ;
		END PORT
	END pin_937
	PIN pin_938
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.17729083665303 0 70.42729083665303 0.25 ;
		END PORT
	END pin_938
	PIN pin_939
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 70.49701195219087 0 70.74701195219087 0.25 ;
		END PORT
	END pin_939
	PIN pin_940
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 70.81673306772872 0 71.06673306772872 0.25 ;
		END PORT
	END pin_940
	PIN pin_941
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 71.13645418326657 0 71.38645418326657 0.25 ;
		END PORT
	END pin_941
	PIN pin_942
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 71.45617529880441 0 71.70617529880441 0.25 ;
		END PORT
	END pin_942
	PIN pin_943
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 71.77589641434226 0 72.02589641434226 0.25 ;
		END PORT
	END pin_943
	PIN pin_944
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 72.0956175298801 0 72.3456175298801 0.25 ;
		END PORT
	END pin_944
	PIN pin_945
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 72.41533864541795 0 72.66533864541795 0.25 ;
		END PORT
	END pin_945
	PIN pin_946
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 72.73505976095579 0 72.98505976095579 0.25 ;
		END PORT
	END pin_946
	PIN pin_947
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 73.05478087649364 0 73.30478087649364 0.25 ;
		END PORT
	END pin_947
	PIN pin_948
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 73.37450199203148 0 73.62450199203148 0.25 ;
		END PORT
	END pin_948
	PIN pin_949
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 73.69422310756933 0 73.94422310756933 0.25 ;
		END PORT
	END pin_949
	PIN pin_950
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.01394422310717 0 74.26394422310717 0.25 ;
		END PORT
	END pin_950
	PIN pin_951
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 74.33366533864502 0 74.58366533864502 0.25 ;
		END PORT
	END pin_951
	PIN pin_952
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 74.65338645418286 0 74.90338645418286 0.25 ;
		END PORT
	END pin_952
	PIN pin_953
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 74.97310756972071 0 75.22310756972071 0.25 ;
		END PORT
	END pin_953
	PIN pin_954
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.29282868525856 0 75.54282868525856 0.25 ;
		END PORT
	END pin_954
	PIN pin_955
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 75.6125498007964 0 75.8625498007964 0.25 ;
		END PORT
	END pin_955
	PIN pin_956
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 75.93227091633425 0 76.18227091633425 0.25 ;
		END PORT
	END pin_956
	PIN pin_957
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 76.25199203187209 0 76.50199203187209 0.25 ;
		END PORT
	END pin_957
	PIN pin_958
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 76.57171314740994 0 76.82171314740994 0.25 ;
		END PORT
	END pin_958
	PIN pin_959
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 76.89143426294778 0 77.14143426294778 0.25 ;
		END PORT
	END pin_959
	PIN pin_960
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 77.21115537848563 0 77.46115537848563 0.25 ;
		END PORT
	END pin_960
	PIN pin_961
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 77.53087649402347 0 77.78087649402347 0.25 ;
		END PORT
	END pin_961
	PIN pin_962
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 77.85059760956132 0 78.10059760956132 0.25 ;
		END PORT
	END pin_962
	PIN pin_963
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 78.17031872509916 0 78.42031872509916 0.25 ;
		END PORT
	END pin_963
	PIN pin_964
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 78.49003984063701 0 78.74003984063701 0.25 ;
		END PORT
	END pin_964
	PIN pin_965
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 78.80976095617486 0 79.05976095617486 0.25 ;
		END PORT
	END pin_965
	PIN pin_966
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.1294820717127 0 79.3794820717127 0.25 ;
		END PORT
	END pin_966
	PIN pin_967
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 79.44920318725055 0 79.69920318725055 0.25 ;
		END PORT
	END pin_967
	PIN pin_968
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 79.76892430278839 0 80.01892430278839 0.25 ;
		END PORT
	END pin_968
	PIN pin_969
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.08864541832624 0 80.33864541832624 0.25 ;
		END PORT
	END pin_969
	PIN pin_970
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.40836653386408 0 80.65836653386408 0.25 ;
		END PORT
	END pin_970
	PIN pin_971
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 80.72808764940193 0 80.97808764940193 0.25 ;
		END PORT
	END pin_971
	PIN pin_972
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 81.04780876493977 0 81.29780876493977 0.25 ;
		END PORT
	END pin_972
	PIN pin_973
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 81.36752988047762 0 81.61752988047762 0.25 ;
		END PORT
	END pin_973
	PIN pin_974
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 81.68725099601546 0 81.93725099601546 0.25 ;
		END PORT
	END pin_974
	PIN pin_975
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.00697211155331 0 82.25697211155331 0.25 ;
		END PORT
	END pin_975
	PIN pin_976
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.32669322709116 0 82.57669322709116 0.25 ;
		END PORT
	END pin_976
	PIN pin_977
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 82.646414342629 0 82.896414342629 0.25 ;
		END PORT
	END pin_977
	PIN pin_978
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 82.96613545816685 0 83.21613545816685 0.25 ;
		END PORT
	END pin_978
	PIN pin_979
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.28585657370469 0 83.53585657370469 0.25 ;
		END PORT
	END pin_979
	PIN pin_980
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 83.60557768924254 0 83.85557768924254 0.25 ;
		END PORT
	END pin_980
	PIN pin_981
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 83.92529880478038 0 84.17529880478038 0.25 ;
		END PORT
	END pin_981
	PIN pin_982
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 84.24501992031823 0 84.49501992031823 0.25 ;
		END PORT
	END pin_982
	PIN pin_983
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 84.56474103585607 0 84.81474103585607 0.25 ;
		END PORT
	END pin_983
	PIN pin_984
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 84.88446215139392 0 85.13446215139392 0.25 ;
		END PORT
	END pin_984
	PIN pin_985
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.20418326693176 0 85.45418326693176 0.25 ;
		END PORT
	END pin_985
	PIN pin_986
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.52390438246961 0 85.77390438246961 0.25 ;
		END PORT
	END pin_986
	PIN pin_987
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 85.84362549800746 0 86.09362549800746 0.25 ;
		END PORT
	END pin_987
	PIN pin_988
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 86.1633466135453 0 86.4133466135453 0.25 ;
		END PORT
	END pin_988
	PIN pin_989
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 86.48306772908315 0 86.73306772908315 0.25 ;
		END PORT
	END pin_989
	PIN pin_990
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 86.80278884462099 0 87.05278884462099 0.25 ;
		END PORT
	END pin_990
	PIN pin_991
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 87.12250996015884 0 87.37250996015884 0.25 ;
		END PORT
	END pin_991
	PIN pin_992
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 87.44223107569668 0 87.69223107569668 0.25 ;
		END PORT
	END pin_992
	PIN pin_993
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 87.76195219123453 0 88.01195219123453 0.25 ;
		END PORT
	END pin_993
	PIN pin_994
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 88.08167330677237 0 88.33167330677237 0.25 ;
		END PORT
	END pin_994
	PIN pin_995
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 88.40139442231022 0 88.65139442231022 0.25 ;
		END PORT
	END pin_995
	PIN pin_996
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 88.72111553784806 0 88.97111553784806 0.25 ;
		END PORT
	END pin_996
	PIN pin_997
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 89.04083665338591 0 89.29083665338591 0.25 ;
		END PORT
	END pin_997
	PIN pin_998
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 89.36055776892375 0 89.61055776892375 0.25 ;
		END PORT
	END pin_998
	PIN pin_999
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 89.6802788844616 0 89.9302788844616 0.25 ;
		END PORT
	END pin_999
END MACRO