MACRO cell_0
	SIZE 100 BY 100 ;
	PIN pin_0
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 63.0 1 64.0 ;
		END PORT
	END pin_0
	PIN pin_1
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 0 36.0 1 37.0 ;
		END PORT
	END pin_1
	PIN pin_2
		DIRECTION OUTPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99 36.0 100 37.0 ;
		END PORT
	END pin_2
	PIN pin_3
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 99 63.0 100 64.0 ;
		END PORT
	END pin_3
	PIN pin_4
		DIRECTION OUTPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 63.0 99 64.0 100 ;
		END PORT
	END pin_4
	PIN pin_5
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 36.0 99 37.0 100 ;
		END PORT
	END pin_5
	PIN pin_6
		DIRECTION INPUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 36.0 0 37.0 1 ;
		END PORT
	END pin_6
	PIN pin_7
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 63.0 0 64.0 1 ;
		END PORT
	END pin_7
END MACRO