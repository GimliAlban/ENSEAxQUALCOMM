MACRO cell_0
	SIZE 100 BY 100 ;
	PIN pin_0
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 0 49.5 1 50.5 ;
		END PORT
	END pin_0
	PIN pin_1
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 99 49.5 100 50.5 ;
		END PORT
	END pin_1
	PIN pin_2
		DIRECTION INPUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 49.5 99 50.5 100 ;
		END PORT
	END pin_2
	PIN pin_3
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 49.5 0 50.5 1 ;
		END PORT
	END pin_3
END MACRO